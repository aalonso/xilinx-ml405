XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���s�J	]ȵ.+�I�uf��`Z�_�~�&�D�R��
$_��;-�Qӈr,���(��	���ĺ--A�Sp��O��emT4����e��h�UDbF_rA�);�Nc5���i�4Ͷ�J4�v�UzX�l���7��}4Uy�@*m���_�rJ�F��9<t��&�O���m �P:M}D!��I
���� ҂d'�}p�n�K���S��5V���(j_������mX ˯��#����F�I�Ǝr�����*��X|�Q'a|����8"�FL7�"�X~�$B�v���UU*4h.�ǃ�c% v;��.41��9v7%6؟��n�qlu#���SQ��{_s\�p�p݉� �t~"�%��̀}��CF ������UT��mZ`�j)�bͅ�$�;��]�G����\��å�x�ӆ���]���ɕmy�����(�v���I��*��5��� a�Ro�Q�G�Q��(��J�9����0�n�6�W$����j�G�&�C}x����lO*���=n�G1��Qo,�2�1�u4��B�ь��7t󻂅��˰���)���/q���vj�$Q��� �9�Fq�a��Pub���Z�������l�P��F*m���+!C1=tp�����)���7�Y�\�7+�8{^��qu�i��![{;TC�}�:����ǯ%�?]t�&=��f/=:f�h�5����a���{�(p�p�5�/		J�g�m��e��FN�Y���XlxVHYEB    1eda     880�NW�Ԓ!x�3��Ts�k�.P�f�����ɹ���YDS���i��-��V�����@-=�B+c�n&H\�Hs�ֻQl�_�IGY�|~�{Hû}�v�Zkiu�d��e�|z |i�R
!2K�Gi�֒��x�K@���q�Ir{j�-��1�X�:?jp[��0P���Ӂ�X�M�ǔ��^1*7v�j���9SJM�A�0���DEJ����t}��%
�9�E��T7DT�)�V��-��<�b�5��z}�I�s�o���ٵ����	���X�p}��F���-��7��쫭c�9���������4g\5+Ʃ�
4�ߴ� ٸ��;�[iEje�jA�+������U������^r�`,F��gET$�k�7IO�r&��ʣx��lLf�S��U"�y���ii��x_�Q����JI\z�l�����a��jH�J6��P��
�����oXs�9�-ue�v2�ï�O0ń{P-��.�8���E���+��
R�&u�O%\��*�q�����y�>߳b2�H���v��OU��-�9�|�f:R��n�
'�E��a/���(�ȩi�yLn�7i6)B�k;[�;��|�9T**Ǣ6��5�����<�c���Q �Vyf�F�]��\�gA2�
��8�S�rO�y��Q��,:Ɣ0Ƿ��[N�c�b���@56�ӢY�D?�n0����:�7l����-K������z�)s�Q���j���!����Jc�K���9�"f��a:��VN������CګKF��L��7�2�ұ:���w�S���-��M`1�\%�A���6�:�L��v��G�ޭ�xTF���*��y=��:��{YD�I����j�i�9�YΧ��bAJ��I����P���֦J���\Nr^ceI1�BhG/Khޤ���[�Z�s���wb�%h
f��,�7;���	d�ms��A��W�����$�<�q4�	ߖ�]��Xl�ؔ�f��$��� ��cA� ��y�I�`�x�T�
���zut�
���2�]�P�Ok�u;�	A
��۴ͼ��?���~��W��S{�5//���	�Mw�o����>�N�7�u��ؤ��Κ�$�n'�:��(�Q3.f�;(�8|�֑��N����5�7ݣP[��T��C#ٱ�̦�
�I;�.ʦ*=��c	fBw�ٜ�:�^�A�Cyq
��2'��-�?�?6P$����xm�&Y���m�2�[��n����9'p�%���6�����:#̎kR�	��u�w�Y@�=ߩ���l+�1�b}�� �'�,�ؽ��T�׫��&%���G���J��a�}�S�$�k�2��8V�OdBi��,�)�oL\ܷo���qu�bf!.D��m7/�.9���HZgX:��G��PpㅃŦ����登�RD4d��[,����a�#y?�SB�f������K��}RT����JH��,���?A�ԙ
����D��1�՜'��b�:�[z1�UaOe�;G\Vާ�1��){��݀����+�ن�|q?I8�8̡��?���w_�G���r4�N8������48q����q����	��Ѐ���˃;���C&h]`R��]�t�K�{��qR X�Cx�I�>�N���)�{��tJ��<���'sO����R�-���M\W�1(��8��F3�dP1�PN�6�(����W@A��H!$�����{��Qb��RBh:�������(�eR��U��+����9�W��Q̳����Avf#|ϳ�Z��m��V�6y%�����pԖ�sbP&��,w\�����c�ٞѪ=�ư����X���N^��rT�Lׅ0�9T	G)G�>�+���-(
cf�D-�;�om|�h.����>ȅP� �#u������1#x��aj^t��/�#��"��@��O�'��#L�A�]�:��_
U�p�#�e?����4@�\������B,��1	s�ʔU����.1E������R�T���נ!�|�E�c��~@,v�����k�?k��b�w7V>;�XA���;3��mS������Ϝo(c����"5���6�{�����]�1�\�.�s��̉\B�p=Lk�E)d8��#n��J�t�