XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���3��2f�rmrհG-��B��c��Ԟ��@B���Jo�W�s�L�M�Nķm�S�j{5�䩬o�]�O���쁈^l�Y�"$���+�I�3AW"<��zM�i���^*��Y���M5�hr�s�tG�� ;��ًp����'N�6y��S-5G��Q��G7Z�'��C��/P��!3B�?�"`>A����xȟ�݂�E [9�����_�pin"u�x��c�?�捈Ѝ	w)�_3�)��e���ש:ڒ�5���Y���c%���X��xsB�}@U��k�����)1��`�\����=�Xڇr�h�\q\x�¶�/e���
�����\wb��wK�t���B�9�+Q�jG6� �|�S��йAEh�k�/\��Pʆ��<|��hd���JeC{�ώ$��Ǣe�@Z���%zTVC���V.���H�SS��H���W�4���j�K����$萑�!����s\j�zR�&�Y����������č�l �a2�s�V���_��h�2�@)T���]N(x�vzOb�V�~�U�\ ��zC�W�C����)>���z˪X�����\!:m4����ǡ���s���Ap��	4�6�`��~������>�T{�C�S��'��Q�j1��"3��ܳN $�p��%\���	)��ه�bFWygݞ��x�Xn�ݦ�lu{�پ7о	��0Ð@(�fڑ8B��Y��+<.�t��-)Nm��L��JRC��NR�L�XlxVHYEB    1e12     920�n!�*׃��ЩY����8����M��N�������~v��Kg$�`�t�0��"������p����cNSb�cU?���D�Æ3d���oa1�� �5�/���5�q́�з�f����򉀽��HpnX?%t�����)4x6�k���?��#�PVc���ؖ���չ���&�h<�e�(ۂ�\�-���B���r�^jܝZH�]9U�Yz�Y�	a�g�E����_�5�o�e�;Ӥg]ˊ
w"��F���jW+!��M���~�>09��י5ϮXV������>��5�Ȳ�ӏ�so*�n2�u@�:{F���יOHf�j9���B2��M���KQ��:�b�L�
l	�����k.#2�a:�O`�!�I]�>�jeg�)k���T)��1�p��o�V`Z�i*�|V���NzG)�FH3�����Ep&M���h�9 �A>���kp����;��� Q`�੄�pr��R.�6��6���Ǹ ��&�"�ϴQ&e����15���,dn�`y�V�d�)�C1��GD%8�*��rK�����U�Wip�q�|W�)�(E��_�������Tչ��Y'po��
��yW!2�A�>�۳@�������o����h*��U��%�� ^��rp�߯�l�ĥ��D#r� ��iE؆���b�@ ����f2:��_����t\�G�6 ^񶨽�|^��3n6��N#N�=ĭC��J7$�����c�I�P;�����]B�*���-Z�l�O��z�V;f�%�JJ=`^���	����B}S��E����J }(�a5[��[�K�Fi5�jK��ʦP�o���܄�>�E"�[��h���3�:J��v"@ѱ6 hfԜ�N"� �=��$�"�V������V�ױh��M�mT�Z?��۟�9�}wA!-Z�v�u��а6E�xN�TN?�y�	����\�����EL�o7�,*�n	j.��j����,�b��:���6�@f�m�%�\���>I��-�/:������sg� ��P%	0zF�{�"��5�@��xt=�w6�R��W���,�k�v��]��3aöFnC��Χ�*�׸^V[I�X��Ss8��Z�}���l�X`�mE�'9^Q_y��@j�$(��_쉑��P8O�>�k�Ɏ�^�,u���h��D�R6>|�(�m!�kΔߕ˃�O�T�%_I�f�%�z�M�S�a��YL;���1���������c�Ek��(��A�+c�3���B_� Z
<�m3��M�Ϯh�޸�Jb��E��sg�����z܂��rE�B������}�	�Ҥ���;9��ʱ��0)�AɡD�!�ő`{��Y���m�����x��Ǻ˄<�GU��"w�wrS�ld�*�<#��3Zə�2t�UrS��;�������G$���X��� ��!E\͠�jR�wR�fhx�'JQ����o�jd���%��T%�aע/�b\>�4SÌ 9#��h�'�d�_[�_4&�!3:f��ua��2B �[k�ċ";˵X[M��d83���������f��?�s��ģ�"Pƺ�.�!�������E`���6�_�l�����!^�S�q5ro�܇{Y��)�ZK~��O�)~w���k��<�&L�+ѥ�f��͢�']��(sd�)q0���޴�f����YDr�o:ɍ���C���`q�Ź�)�Vڧ���� ����Q���^����o�eR?ܰ�ܺ����a�(ȴlt�����X�DG.�5�i�c�s�n�i� .*�o��`�x+u�k3��������<��iC��Q� �j�1%*t���,�S�R8�i���!K��}g(��6�!"=P��;
d���K�Gi���z/l�'�_�/Xj\H�gi��>`�Ø%�r�uQ�ܵ�ד�.v���K]I7��&9�к�|n����d��'U��S��BR}���b�T�f�](���7�ʗi�?ϝJ�x��/E�=�M6>����G</:�*��[�]��|F?�8�N��N�K�H��}ԲÿYlJ'���ի�zCRZ����k;���^Y٫#�-��y��ݪkwr٭`A�6�Vy���h�!�1n>�p�B6�� �*���� �J��m�����h`��Ah*����8�n�^h���b����Q�� `������$B�2��ũ���r0�F���[�5���sJ��^(�P�*b���bJ���������:���H��O{�Q���y�&��P��Òꬒ�LS���@���S�? Z�_�D�