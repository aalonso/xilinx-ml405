XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����m'�|?���n�uqB�;�HF��H�x��#;�;��<�V>z�!�ة��q���Z����l[�����{�����8���9Q�u�\#X��A��"9����Eo��O�&V=XΦ�T�������W�` �SYu�
L����U�9벻(��>q��$������o�/�ּ�R��~��2���rh$�,1]zН�4�si+&�X�*��sP�~���?ϬҎ���+�K��H:d��c� ��������K���1=_/��a���>T�;�ũ�~;�s{�P��<?�{�A���T�0�!��{�ʘ+�_��_$�Cݕ�9�(:�� ��P�-j��X+c��t7�`,�A���c���+v0ie[�W}�Àjũ��u�ID����:b�=%�-����,-�yI/(�\=yv+X�@��%/���� ם�v�%��:�F��[�x�1�� o�� �69"x>9� ��(8MR�#�j�:��_W�A� >��-B5�yc'�RH�M��0=<3��T7��U�&�+�����Fa8�R*��+��-aP�������]�[Gs�v���~���DYnI\�#��N g~���1OF,ǻ���Q��=��1m �J��xW{�JF{�.�0��җ�=&�ca=��&���ĺ�^Yc���3%	�b��z݃JTl�SlArqп1�a���=����'����₁�Wk�/���V%%�L�L�UȨI�c@�����/"`��0lO�*��&XlxVHYEB    bd1a    1920%�4� �e�ά����L+|�#;!y|��8���@Ob�����uY�����C�=��.ee�8:e�j�g�h>��\]��3 ��~�IM���_Ѓ��՘�z�K���`��3��Vο~���ǃ�
�*�`��3\�Y=�f��/�Jh��F�Z�z�3֮��(����'a�0v3f5�9����_T
>p��O��ܽ�L�w�"���1�-Lp�b����1�n'鱄o�,�x[�JL�
Y\�
n�����0Q�!3����^��_�}-��;�����ug��nnb��Y��rg'\�/�@�a�î�s�~�z��(��2��� n�OQ���ꛩ���pO��ᆭ�ς�]r$*D�u��Hx��r/�/V�W�jz(�{�ٓ� ���w7�-�����.�����Bs�"��5�K$T�I�^Ѥ�e�.�����3�Ӑ�[(y�֚�xxy�Ex�MG�/��������6�A��҆��X����?&O��о?�6'�Q���/�.�zic�/j�K�c!)�b�F��l�O_����\���MV5�p��.z�p��QK�l��waa���&�^O�G��%r�q�gwБ�BR7ڧ[V���0� �k(�
7�w�uA�S�ϡ"vs�x�ݻ�W��FV[���_n���0��0�t�MA"��-�t����'
���qYn��y�g�- 7i6ӧax�؞���Y�\�V�̦���xt'����F�G?p�7�|�}���R��!S}�?-5��e�����7�6�ys�ϠUoʉ�'�h|`�����t�}!/	`��[�X������Tw�/'�߈́k�� Z�Q��˅@AC�6�*0�־�A�B�X�QFٽ"b+7�ovG�:f�B6G��~��⁶�z>�+˅��<�_0����?zy��a=Ͳ.;q���r�=��Z�o�AqQ�N;�c@m#-��BY�`i�(f���'�PRs\쎔eMe{�����xL�x^�S�%���D� X-���o} �%;�ƨ��&�:_^�sZѵP����p��ճXh��Uͳ�1��5}��emt�1����_�!�W�
�XT{�z��.d�KQH_�Nq*;�v�LBu��%D���꥿<9]�$��P�9.=:���v�G o�+[ϒd^t��THֵ*�X��uq_B�?�t���8�,�D�ޏ�~G�~=�T���Qg\�^^^�؁�'���lŏ�Ad=(��Zsas��v��~n�T	�_^c,��C �nAۊ���^vd�a^� Xɽ&:�� �k��|�7zW��b�zgsf�II�j` �Ӥ`�ׄs�!����Ej���3�CxЖ�����`���p3�/s?'� �"=>�1��C���?��N���Eתo	�Gp@�����Hθ{���/�"{=�٣�J�1�Sx+KF�Q�EH�'?�����9"WڙK�is"���z �Wp����#	ۢ�����g���/��s����4ɫ��?S_�6�)@u }CS ����Z�28����ع����#P�vcY�K���W�[0��+3�T,[��oT�㨌�P�ը�G��|����Ve�����Od�O%�r {��7�a�*$��U���~T����R��X^��d�YE�7�m�m��	��cJ���+81T?CI���hk��ݵWPT�=)��A3���j�q3���R@�_��;��� �jm�Gx��XW��<%�?��H�M{��d2�46��h������{�+]�b���[S���ryr"Zua���*���T�K��m�:�'^�C��$,/6FX�-�l����V���3C'%�\en2Y��l^�J�d��"���C�u`$�*�1_$��K����qs.1���F˂{�]�9_#f�@�����AK8XSs%j��l5�İl����t^g�_���PgF]4dH����~�k��Z(%?��T�Ȩ��A�:�ڪ��IsQwہ��x��v%���*�
?�����5ȣ�x�eA��� ��.a�"XA�`X��.���nqnx�):�Θm%�4���֟�)�6o��^�y��%���5�b���|@��h�?୊����Β�:�sN�[8i�G&��rs`����bp ��5�F�Ip�q})�'hx�l��?Ej��B���C�f-�����LW]��\�����	�Βj�����х�~�,�PD	��<~l������=�%:ӇXʊ>"��8�p'�4��x^ ���N�@�6��������u���8�ZE�K~�l\�Z��;�~ǣR��N��-���P��_I�	g� ��s�049)7����eJ֙E?��[ʝ�j���Iޚs���������[f���5Һ��8o�׋�'Sa�%YѠ�th�oz�}/p_'<��R�����fn>��$ކ��?B2�A�����e���x㐃#m`�/��b4����f������%$n�c`��B�'�2���Q.$��<qH}[�)��!�< Ô��ǋKm�˃HG���P;�����w�ko.��^�6C�qOYٹ��=�ט��<\�<v�C��7��9PBK���ߍ?X�1��*B��Z:��}ՏU���H�W������S!��:��( ���J�5BF�$�z{���pzh��L'��������g���n�D�P[Ǖz�zO�I%�����_�������L��~ ֨,�� ����p7.����.�աt�����~��֥��}*�R1���[�g��b%��9��\3�V�ڝ�Evai���/3Gf��{�1�o�F*�+n�A�d���$�嚎�׬$�<^�_�r����_Ld�R�y��N�(z�4��r�����mܦ|yM"w�x�a�%�,Ǣ_�X���F�
Nm'��.��Pc�ӫq��g��2�њ��nt6���>�*'q��{%��7 � C�z|�TsR)��>�ן���������ց��Su����r?/M]��&���G*��m���ؔ#>=jb�`V�K��_{jʎ�}g��;w4�>�0�&�[\T-��{��4���9�=f��ߪ6;g���!V j�H���_-�$��C�%�Ko��gP�I�v�Ǥ�ۮ��ꪷ�[����7�F����W�'
���&�>i]g!�bj���t_�c�^qέh����/R¬�����~Y�:��L���e��?����A�C��BE0����������n��7�UU� R�*�s�|�L��**�����~�K�����^`\|L�gP+Na��F}��M]^�u�͜.-�A��{F)�o�j��5���V1 �d����Ħfz�(��^B��П��,d��>���)F�̂��A�)����R[Db��R��(�c�Ax���Q,e��ޚ�=�D��C1� ��#`�C����.�S@֌�˃���>�`4U���=�7�ȁ��*�7?/��2�
��@�U�jr�����}Pi>D�Id�H��<��Fg�]�[*��0�_�z�m�Q"�<�t���]��?�	�n+�H��?}����VoTX~³�d_���S�(��YddG7���ʾ"��ı�&+AT�·l�O,e@e0�|��h4b�r=v�Dxz��^�m����i���$%�/7�C.��擴�5T���eV�͗;]Ǯc��y�}L�9d�u�Q91��t�O��s� �~byXF�a�ﶆ��u��\�	$��
�	�-��;a���>r�P�́������r��`ߪ��8�/ڗj�SC��π�^2��D�A�aF��&o�P#QEr|��bKR��S��c �%��&KM�&��4�@[�ur��+W�j�30_9�w��4@�S�>qk��讃�,)����8/����|�yd�i��{P_���y���/�#�*�*�DE�L板�]�4�F[�G#T}�7-���/��a����*d��>$>��_hːYJ%�u��s}0�t:�"g�ļ�=:�D�:uH잩F��e�8����E����y#�j܋��M�U��iz�������I���wX��Z�{�3��Ȱ���C%q@C��l�SXkL;-='Rvu�E�gt��X����ю��[���e,�VEUU���㰵oYZ�����3��]����=��z�v`i�'J;h���l����XIA9je�2_6��>H�Fk�)�N/O�� ����xW���!	�����7�z�=
�d���\'r��B�?R�4�p'�l�(���j���%� ��B�]��{���j���%�G2�}n��Z3QG5j��nu��0\x�_�7h��kw+d�����6������������Ņ2�WMD��3zp!y}�o���'���5�+��_{.JI�Bĸ��T����i�$�B���ػ5��[�9 ."2{�޹:���;��B�R���E��g�������m�/�ȶ�]�����[�@�W���f��@S��(������T�y��D���R5ak �"�������Z�N�v{*�9�5D2�7~� �D.J��4ɦ�z��HO�V�b�Zs�|+zbgo"+%��ϩ��G���l�����=;�'m�=�+���SnC�ArN_t�'\|�@�s��\� ��b�|5�u�}ӷ!IL�;r�7%g��x���h����݇�tV�2�PG��<1/3��1ͬ���n�3�2�@aJ^�<�{���j��A��^�a���X򡹴SߟN��+�1�KbY���P��}�m����p�ɒmR�"m#P/�.��uD�b�첏�T�q�}reI��������3������w-���K��:�~M28ɟ�^� ��2�MI�)�n�|<�j>.�M�jJB����ݛ~������*�mm�C���iR��0T���H�E�2Dq�/�@*+E!����S'A6�r3S�ai��ү��˙�]�{����W&"��i �ZK�	m8�N�����\4d+7�+7+�8�ĳa�3�ެ ��w��;���]:b}ۺ����p�>��K�:Bc�p��O
{i��w�&��Ǫrj�Ng[_^�!�W(ȅ�ʑU rK>B,�wU��ֲ��*�M
K���d�`q^�P���x{��BM�h�m�*}���N�54)۔���t���G�s�ܜ��XQh.wX��k���}Y�q��mt�z.j�x׏�	�C�'Ɲ�50��J��Ӿ6t�.^I�:f�i��xi _;C���;�_e��rno��IMJH�h��zO��5ĝ}�L�d�!�Sv�M�r}��6ėk	�\CK�ĪnV�U��BC��f&^�S{wvt�1�^j��T�yJ�E7�[qΤ�̭`D||���ҳXS�Zr�ƨ�w�o%_���H�Q�I�y0fm����f�\dl9�d��?��a�o3 sAu���0������;�f�x��J�� ����K�I:,����g`��o[�ωѣ6w�j��ػ�sN�ϑI6���_?�������N���^�$b���s��>�A7�������u��l��-�����������j�m��pn��f���Z�k�3���t��jS���`G��d�`�-k�bgV:X����*�y�j8F��Gi�x���-L�Ӳ?k�LDnkk8���S��>�%t	J�>W�'<�d�t��OL�� �[��N�����Σt���S��$
�!�VQ@)ڴ ��%�(N�_��p��`�ƭ��{�%�x��TlL�p�
Ý����k����a>�?����`g��w)nC/�D8\.�����PfXLTp�`�'�0���{��5K��㟸b b���{n5�;��;�NƓ�'���awi/J���4w���#� 2�mp���R_�n�"���Ö�C�u"���NE�����|41���J�T����.U_5���&*->'�g��2ΏA�"V�5��պ� ��z�X��CP<f��,����d�a����P���O��ӤN�}�c�ڏ�-�$Ze�����g͓�;o��Gy�w�f\�$��4d�:��n��:j�
"zy�����#�H���C9��Y�	"�{�ێQg�(�e�5�����Q�	�2��z��ȧ+�Ʌ	9z͑_K�b�/n�KߩL��2L�#��X��B�� ٠�n,�K�W�P�%�� O^e��������vc��&�N�d���ۋF�p;���U����$<�UpkP���3���M7��6���5�80VĂm��d���0Ж���X3OZ��'��~s�Ut2�z2gzkJ����.���q	���Cj���Ar�d�L�=9>��b$џ��!���?��@�KD��S�Q\��[��s
*�.�
��'y���,��Mj+��u��yL.�r׃S����Z�3�