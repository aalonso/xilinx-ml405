XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ճ�m�r	�a 8Av�բ���B��Ul0~$*���7�7����%���pr��i�قi����<T�Mx���3��3��T�p�"m3"[K�짭�ްޮJ�M�U����\����]L����O���z���Yx<�hL��M.��X�3�ϞZ�ܪ�T���M[�	Nz ��=d9��*Cg��E����%.6��Йj�.�S?�v<��˴�Zu�T��$H����e�4*��./3�""^�>���q$%�����V���ue����f1�,Bkm��v��W5���n�,����.D�D��z�\-� O�#��rN=��[wh��p^ zÿw[IeK��n�zlٲ3��dIc!�	��Rϗ���`�c�v�-�_~0�Lh
�`-a�[ܾ�3�7mm�E���.�Y�ڈb���lAv�
h}�U$u�^�\��t��U���T )�)L1�JT�>� @ٜڵs���c���΄L��a�����)q�Z2�_��P���#C],�w����:l���s��J=}��*��h�T9��ÿ׍�Ri��Q1���}3��# ��H^u��r.YZ)S�J}Sr�Lb:���gXU��L��9���O���7%�����n?)�2��}���R��� ��!�Q�����u!�C7s-����,8�E�Ё���SdR\ܲiX"����M+�/+܇��C�a=�:�C�>@�V��̈�]����Xj�ҏ�l:5������GjSHR@e3W�oXlxVHYEB    fa00    2620�,�6��+AbT��2۴7��Bdb�KҩG8I-K���"X��}l.�/��Q�J9����Tyn²�X�}hK	�B�--�u�c6Zqq��r��F;�� ���QW����Oy��p���&���'�S��{Ћ�ݘ�a̸���s�'��1�R�&ÀolH�Pe'Hz�����<��(]��+ࡀ4�UY˟דA�9R��5E��V��F2��K���JI�`����e*I7V�+��uc�y|���+>e�i���W�Xy���}˽�r'�� ���.�=^�j�PK"���#����D�C���U�d�L/U�h� ��,イ����p��Vzb��� .�㒔p�i9�(��ʲ_.��ԫuw�1hQ��W4�Sx@�ϒ(Y�m��mcj�ٞ�z7O�ʹ�О����F��na����|�h���RSE��	.���0��n�ག�ĉƷ������=-j�ɮ�Ll=���$N)R�����R]�ߜ�¸��0����)��A�D������Q]��:R�0<aTd/`B8�P�o&R���Z�ϧLR�'�L����aW�����`��)���pz@�5���j���XS}ɼ8�s�N�-܁>+�Q2L��ܞ�ER(LU"�n�{yv�a�C$��S��^�T}���ψ;FR�#��F�`3�I�����e�P�pLD$�`�R�	W9�G�0%�'�x�X��Gy
�Wu�;��B��y��l��\�+�TU��7�8�����r�O'Ϛ�C�V�{��Xݰa�Zʹ ĄG��%Ƭ�e�,V��YT�2H�9	�憙׉����	j	�Wݼ���%�|q[�x٣��
���A��I�����P:�A�i/=�|b$�%���ԄrI�����+�/^�g���vU䊮�ꉂ��,��tn��pK%]n������`܋^"[�+U��ܡX�Tǎ~⃇��l0��
���A<���uM�l�t"�^��M��<j|2��Vu��N��*��A�j�f��K5� �:�ݾ�r?�[���ޡGqgyf����NYH �+�J��OD�ٗ��'�]W��N��(6EoS�����.J�2��/� ��Ԡgv��g�q��1Y�\;;9�"����+��W3K�����#���6�aPR�h�@�`��ވ8�vtX��r$�5�}7i�E��q�D��s��L� Թ*o.���=�>q��}ۇ{�����a�r�C�͂w�wg�|�qW\��.C+[�x���y���*��c{�L��e��9�V����4wN�"P�y�َ�C'���gI���`�����`$�;�1T��e�z^397W҂�u�0`�A_C�A���9����#�X�>�`'�1-/3#����ܝ��b�PQ�O�嘏n��+-E�h@��z�j������K>)Z�A0'�47���R�� Z~��I���k*q�ۻ|�v����chR���+��.J�-{m�-����"=��g��e��s��Ҫ�u�ʥ�������=f#^9Q�ƹ�=Y�W�~�hh�2 y��	p�ϷR����#ިYZKʀ��/��P�U�X���72��a#�����b^�G�{v�{K��M�l�^�bԓ��������"��/]O�'٬����m�#��!!�н�LZyC<ON�$��c�G�o��R��|�=��L��L���^9?��Z�����~�ܢr���0I�+S�G�,�Z�{�����õ_�V��r��p>,#*+C�b��]����"����Uq�Mq=�:������=�8��OF~�g��w�k���u��f��^ ���)���+{��~� 7!W?�<�J_�?�[�����_���;cDk�PL�i�cJ�&L�U�dН����v/ͬ)�W�.�2��Dt�^+$�����2-ȷ_���Ԯ?�G��X3�gb������K���l�n�={xl�?�c�!v��I��;���l��E����r]ő�xX3]����к��T�q��Cǹ}��Τ��59�cM�
�PD	���3A�S��8�����h�]%�ȂV��}�p�Z�l�4�!:���ί�W~��Op�U�H���aAn�#�6Ŕ��ِ8Ȯ��F������n�j��Ԇ�?��o�3ٽ0ڶj�sW�NڪF텆B���@�z~"��j����R��ԒC�2���:�Ѓ��"�ɫ:��6؞f1�S��~ R���۴Pv��v���+"�d��g^Z9�`e��
?�`�H�.�5q_@g&9�1u�S��5�_h�"z��а�S���,Qނ�ˤ(������,���Gd��H�[�	�٩��Z��9�����Iߞ�=-3c)���#��!���Y!eї�f5	�x`*bbxwź,]t�.�MY���c�kۈ�����?7=hw��OC��8l�ű�d�7� Lb*�,�8��'�, ��{@	�SS(�I�����Ŋ>;���/�`k~5��.���I2�����_�ߌ��_���9!���ؼ��M�|�}�J�3g]��A1l�>�Ե��󧿎�P��@��VE��B��u���V��uo��&X�`-{ԧ������`��+/�r;�|�R�}���ږ9��E�2�nM�HPR�OѸ��vҼ���ӽ�z�]����W��D �Y)�	!XLįٓ�;��I�iyZ�b��+)ZK"p�bp��6�5<����0�cߕ�����8~�W БOcJ�����}�����U�}���i5J���?`�_�$��t��ޖ�b�T�e9Jw^����!-"�"q��!�Vb<����vS�g5[���m&�rϟy���.�+��y�
��$�����\�P�ŀ1u�P�(��K*��LdWG����c'��%G/O���Oc�k�t�@���W�h&�� ߄��Q�w-�i�����t a4����0`���"	���>88�)��J�]Cn�I|��Y���H��R�i�I����LV��I�-�J^j~�݀�:0�#� �|�`��Ʀ���r�C	-�Oۥ��g�z&�w���|���|�1kP۶s�?u������I3����&�1�"M�2��3ژx8�jC|5�Q�j��Q�"���Z&h�h �X e�0��95�B�Y��T�3*�-����!C�Q�E�쎞T��i8yP�>cd��.iğVNpZ��	��1+��2K��J���!�����X7�5,cg��}4��w��ݙw�	������pҀ|�ĉ �K��� �������Շ�����+�{���&վe�0�z�ͲV4��������5�E:��/;QZl*�+�#z �^e�h�GLRD J*]t;�h��I�.Mn��Y�m�[��s�5<]�J�Z�4%Vkc����e`W]����]�������
�Z�u�W�B���=Іw�t�m��*a����A1ֆ^�rVd�4z8lR�
3%	�V�w�?��?��ʘ���ln�#f�� 3/�$��hj��v}n�y=S��i;o�qa_��F�`*V�	�ۥ���G�po������>3s�f���Zu��zy��������Y���"�9���P�/��E���`��j���R.�Q�[��l�p�Ce者� Լ$@����(�z�̽2�R*�.؏=�a�
*� z�F��S�$Wk��b���혽܆/CIq�?
��2#*<�[���e�4������7x���8�:+�0}��9c�HJ=���gk�hc��t���[�%ƚ�E�U���DCȞR�w�9�_xt.Ң�0{1��:��Q93������'N���a�S��a��ꁿ6]�H��DS���ճ-
2CB�gL`����1���N�� ~�}���"�&)1Ʒj�K�r�����X v�|$?땓3�o���돢����%m�d�Ona�� 4�t_�*��6uvx`7Q8���su]��'&q�mB������u��K![{��S޼���N�: Nz8s"(�_��l��f�~�Xa���,��H��t�pVM6��o�|0SKx&l��5�G��!�A��}Y����׊�(
�:�x̶>|�W$ jğ& �o�HLb��۝�|�EwG�h�D:��+�R%��n̭
��,z�:����� ���NP�06��".F��!\\�2�q������������3 �@T�#<`��7��?�sE����z�d�dq�7��}�%��"�KAm���2�@y�Yc*�E��ўM��
�RRч��Y�n7�$&QQ���$��g;�k�S����T;�h��>⢜��lAB�;��e������1�bL�����m���5ĕȻVI ɺ=Rbك~,��|C�z��0PRb��i4��I*���i%|��L����_	�$¨�S$��.u�H,�ܪ�ȴ+9�ؠ�����@�2'J�OXt{��N�8���y����|��]�DV��X�ue38�d_G�7������)7����P�Ȅ��Z��M���o�'�z��l',�J1�5Y�D�Y��`y��<��Ꙃ�RLk2`'� ���1nJg�K�nN�{@�/�%:��:�i�zlN	ܚT�DBaď���Y����V�	�h��B�Z&�Ȳ}�Q�t\���>���'�ウq-_A9����rh��l�<3���I���3�îv
���*b�\��,wc���ِ�a�X��4�g7���R�Ԫ�����5�9��~�`�����PO�\[?>W?�
3�6_�`/i�v�b���z��f��9�]ۚ����Xv��捅]u�.]E�U Ȑ�0Z
��E'�|��v"��X}2W��&�p4�p��)���j}���x�<*>70$AEK��3(EPH+�G'rc�:K���(��N�{���F$����T�I�]��k�'��R%`���'�Һ�%��&>�EK�0�G"�T��N��=g���|��kޓܚQ�����/,h"d� Y}\#>����I�E6�݋�M���*�{�]�Fl��B w��ɼ�0�[I�����*���_�5�7��.}�����X˩;u�'p�pCF����f(� �h�.'L��$�V0�Y2����pK�&�%^;o�*y����-q���Gy��n�������$Z�(���-I�S�;>�U���}i�B(��_!�-1	��С�JN��ѝ��KB��� ��	E�U4w����v�ݮ/5�ГrX��n$)��vƭy�}�����.T�I��(/%�O��w�5�n���۔r"G���'�P��YZ3�.�k��moA���*i�z���u��Q��5�s���<��n�	o����3:@yV�':>�� �`ṘF[6�&��h@�5u٩�7?�1vx7.�6�{��`X��A��1�fJ}�>�(��sǨON�M���ͤ�S91ڞs�$�"I�q��S��Lw�sN7���ڌ�	Ҟ�������O��� Ĉ��v2-1�	�'P.x6<��S#�k�j��DxD��K��k͚z�:N���t�~ߏ�\���|�jF�(��%�W"�&�G^xXB���q�y�������쒦�R7Y�n�3��T/T���?�:ɇܲ�O�P�bs�G ��H���%^�;gJ�u�+���6k@un�}�#�jNE����478���6�b3����٣)(W��x��+�泙�|Nk\oO��O@G�Np��ӏr�R��45����WE|"�
�Q������B�^W�f�1!/��[���!1�ŷ��"[D��Ω#�WK�Y� 4W�^��� Kة��D��E��+_R
_?��_Ph@�V�,S@(�j@)�Y�+d�bVw�:�G��g���i�@W7�d���������H��l�*M��� �����������4�.3��{'�����z�x����ՈO;��BϚ'O��6�G�=Ӻ��9�E���D�ZS��F�4��ǧ.��{KZWլ�Y���O�`����򈦆�|E�TΠ扈0=�ܢ@�>�Ȟ�=��{K���4#�L[M䆰�y*´h[�0��R�	DD�>�j����Y6��sh�-R��}�N<�Gݿpn��H�N��w~�Ɨ�/��Eݾ�5o׾yÄ�s�SF�3�5�i�5}�n���9$�
PH
p'�4FuR���yc���l2}H��;췠�؀�D�U����c���R���x���BQߠ�$s鲝�8����"�1�S`�qҀ��O�g_�}�2�����cl7C�0�E����-�B�V���H3����A���o^T�S�Tܚ�ۋJ�ؾ љ�l�\�?��
i:�Xd��B���I ��P�b� O��Ԗ���`�=sk���>����Q�70����Z�{Z�Ŵ`�
/�t��ˉ��@���4�]v�1���Y�(������~	X�W��O:��� �p���G��{��G'��'� ��[���
Cz��Kq$�ݹ�|�O"����8���٠@�3G6i���֓V, ���0��P���:=5�s�`ugEz�ۉN8|�݄j�H�8}�f��u5S׈*,k&?ʊZ~ytQr��j%���������|'�
-_c�齕�ŕ>� sK*&\6Hg��b�u���:��r�3C�����N�TpO�8�لH�6�>´���Ws�սs���יt�����T��Ϸ�A_����=��������z�	96	vQ?��z]�F���멼�ت/��\�;DI�K����mC?JuO�N 6Ժ��T��uw�\��L����KT��P�9��^��N9u>�yFD(e��I4M�Ș�S7$�+�����J�*K2�"t�w~����-��]�0-�4J��udrxU�D@ �cE�%��6�P�vn�����8O6g��A,�J���J�tf̺'�|z ���^���-=�z�Ƃ��-��}�"^���d�(N��3h�٤�'���)������$��|r�j$��l-T��\��ʛ�l!b�,�H��K;�-�t̂;5nx�[��9Ύy�U�d8�S�i�����)���x����	.��k�psn�6�H�OE#\I~t��O�(tE�y圾��W�,[�
~�..�j���Fm,Ԟ����fr��Q9���t��sB���?�A�����7�`o_���-�#�]I�}�t��c�hW�Woh�:��z�Ä�my��Q 4j���dz��/�.~���S�Jj�%OU���U48y-�󺱹�MN!ޒ*o[U�9���,��)].�9��/$2֟)�}�t�q���	Ԓ$X\;���_^��:8����Q�����um���MHo�9G�Yo_΁8sR\2�!���z^s��ֿ���ߪ��i%΂RPu6���O�R	�~C�ӕ�uW{�PU%
A���J9H1B��j
�u8��@.j*}ޓ��r@�QH?��ϻ|��J���z��oў�\E�D1YDsRA3
�_�~���T8]�Drڤ������������ ��gDհ-j��}�-���@�Y*�,�F����7�m�X�S]|��s�K�2#�\�����\G�,����8\y1��9t�	Uw�5eB��#N��NA����(��΁ !6XjI=ٌ�_������c_���~R�:���C�3K���֌'F%�����K�덏Z�V���P�3<��my��
�|m�3������O��q�zf_*زNb�)-R;�A+f��~ϑ!��f������͕k���'$��s.����Ƭk�]�-=-�A�+XS��9�?���|�6��vs������C�/k�-'I�.��w�����H��Ɣ7{~ ��A�陵������|	p��l�oU��.����� �u��qӢ�?H�R8�>Nq��Ù�F�K�$��zؐd�1<
!�Oе�_`�\�K؋h��N��b;վ�h�j�]��x�uV�s܍�ؼ�<*,1d�4-2Ɓ��Ӗk0Zk��a�E�w�Gp6�\��5��o
��T� �7�b�<�v7t��;jh��˱�3!����@��R�ْ�N����e���+�p�&tsGW����줒]!��L-kO�9��x�, ��D�ɤ��gW$-�o�+�ཛྷ]��}�KX�;%�%����4��.m�Oy��hמxk���70G8t5����{�+���Κ*��� ��e:�<��Y��d�~6��EDE��sܵ�Z G�*�����)|��ߞ9
��T$-f�j'�����!�W�ܔ�7�qӝ��ه2�C���Yj�I�H�K���x+x��߶Q�@8��"��qLďW�g`�g{��͌�0���oň�M^C��z�s'��,��(�ZF4����r�9���dg΋�����=���:3�襃�J��ܞ�W��}�W�8��1F�j��{��=��� )�����:9f�9���3�k=��R2��niL�n{̳��s]8I�a��N�}(Zpʕ�r�_�Ԕ�'3��M�;�G�T��\~��ň��1|�����g�ir�
����7����T�w�qX��iuЋ�\�*��E_d�1͏�j��B��?�f�It��^�|O��"�𻗭N,`K���5@S��%�Ú���W ӮC'��m����k�p��1�Z �J����C5�\�_Jݸ����cW��)��&���m%"ύk��bόy�g�G����˧��V�N6������<�>~� ��K�5^�p�FU���G�����s�+�]�h
)�ZNWIj����*�I�]�*@�7�+��fZ2`�dT�۾�\�:�KQ�.��k��N���RA�����Ҩ�;qe<��9��|X
z,١[P�v�6�bq�2����2ؑ��C�5���߼�.��s�´oUmr�_��3����Ej�X����A�%�xv)+g�~����R�E����z���C���ā�%��a�$���f�C:i�_�q�ۤ�;\F �[E�ˊ�r�0d�y��g�;��$XɸeE]h��Θ	���ݰ>m�o|A��1�ҭ�9Z�������� U5�%\(��o���(�Tf��i\)V[J��t�@�f���9Fh�T����7��~����VR{�
14�|3���*t/y�s���HE���^G)���aδ�cy<[������Cn���LBU�;����*�:�0��O�@K?��Ū[�l �W�z^cb|�b	l�����ϛb�2�ua�A�}�:��PL�r�=��Ax9SѼ�jo��S��O���k;M��T�2+x���a��hIeiF�p� P��!��UP�o�'6l��1���,���eʘ����t	ڡ����'��[�pk�LCc���8T�OMq�����cY��Q�A.�#n��\��3>��oRIk׻���g����}<�Bv�h)������*�W(K���	ޤ���z�c+�ib�CwH��X��'�u�)�1S�m<�y5�U�o| ��(
��%'%)���}2�8O������9�)�E�<�Ȱ?Tӱ���xS���Y�w����7�q�d��O�O����������amIsHV��鸼~p'�cVZ���b�w��sL�T
4�b�-(� ʦR�4�f��ݵk̆-�|@�-XlxVHYEB    37e0     ba0�e��\q��ܥ����`����Z��,����'̛|�-c������[0,��c�`s1���>7���'N�9�B�3�������Hw.v��f)����C�׮�{�V���5�L��24d%N����,����uˊBy��nf0 �촢M��fR��Ct�O"L��B�����Ć�YU�nCL�J�.E������]��Y������3��g���eM̉�>�	h�v}��̐�~���t3�'S�)u�t}���ͻ��y���a�o�D!�iߐ���|?
�e|�1���m���<0 σUL%��%�o!<��'�ۤ�(�b��w����\��`���#"��ɀ��PF(ҙG��J ��8��1�3j�3��?�bÔH+3<¹�1�b���@'ݗUFۮ(DBq�8�N,�1��q��o�w�H\Y�9�hY�_����@�Q`����4��^ɰ~[�V�h�1�K��Uҏ�g��<��&Ӳ�^>��߸/�J@B1���ɲ�K��i�d�U���yz�Ш��"ମ��?\�����.��a�,vl0U����fO��e��Y�Ƀ�� >��=�笘�MD�CY]����pRl���d�>
@t�3f��;$6�Y�Hf���0#_����	�:Ȅ��g���a��˖���|0yVG)� �/˹ ��Fޜ�=�	Xm�=Ru�u���%y�),ՠ�'/*��l_���+�hR�	9_��'��~��F-�P���~����l�ю[�t�RIU
ء2R͏!���ի1F'�����O�T� �i�����Yb����	ּ��l�f�J?`F�s�8��ʉ���o�jگ�J��sٍ �ւ=2����fTmד��^�`q���V�!s�}�R�n�1��ЬC�@R����Ӹp��i3Ȳ�a/���w>���s�����&{��\c9�g��Esް�'r�Ѱ�7	��I��c�숏n����=�J� �����Y��1Y�9�^p���n�I�%�L�t�}��@����[�dz��fkZ._���헮}q�Ԝ�eR'ǤW ��æ�U!���w��7r�%���Z����h�rڧ�;�R]�sXjo�g(,�!�$������g ���0��e���ۿ�3�y��3o�
�{jD�jV+��� ��e6G-1��;�Kw���z�u
�M>��~��J(H$�,m����W��s���&��_�zN)�-M�%�ʿ���-����9|��#�@���@Y�'��\���ό�S�vC�m��
��X`M-�ۏ]����ۙ<C�|�9(�J_.ne#�G�5�ך��>��<{��4-�]X��YT�Y	
(U,�-;�B�}���S����O���n�2�g�S��Ð�����R���䅌��(����Wئ���	V1�4�¦�~��b�.���3�<�T]R|�����
�*5�*�`4���~4HyDk2:������ϵɐ��ɀ{�:S�_�dP�A*���R=Z�T{�:@��8wV�T#9i�����n�M_@F]9��J�L����u�ߺF���]���R�MB��/y�E]�4N�6��<i4�I"��]֌���.�t�d/&��=�z��%uww��,l�]WcV �^���d�+�����'�-���T6��N� �Ӟz��\qJ�����mV;�Q�uܢ�4��������k*�|�eYk��m�6M����͘��-J�\��GJ$�8�(��j������»�zR�BZ�Y5Z\"ɽ�|����f �7F��L-#�P����� �rC�"5���I?w��!F�?�7r�2�K�l�p���&s%R��v"�L>^�?���V��r;���3j��T9I:��6����.H�-[C����K�j��PfC�x�1���au��\-�D�Ƚp�,�p*W�.�lv���&��؜�:�K�'�9�M8}�,��C�8��Vf��h�",�m���m��l�����.�xm&�~ P�+˺�_�]3��Rm�z�V@^��J�ѦYC����C����˘A>s�ϴW2��4���v赽揷 ���(��!J��<�݂�r1o�:���}��A���I�fD|�d�+>h`��X�xjvɡ���ur]RW�ǳ���[#1@DM��Yb�
_73eo0�A��C�����7Aٓr��{T��ٻ�����M��gt��[��5�v(	��+~UD���;�`�h�§��x��Ex��.��(�f'���i����<�Y&��&���.�4����w?V�������.A,
V�T��W�B���oHK*���C���F�@�Q���5��:�����ԏ��H��y�Gg�#������Z��5/�X3))�Ż)` h�5��QZ��U_�L��7�]�'�6��	Ą��F�Ne�5����q��}3X���{�oE�������@E_?�{o�&�L�����4�if��zǅR�@V��5�۳"z�N׳���r�J_�����#ty�e��O%��I�SHt/ 
���/�xj�0g��K*�c��P#N٧�]�k���*/�k��g�!�t�NqB'�mNOo6�ꓷ�i�>�s�U�5��C9Ġѝ6�[= ��z�Q#6:)����їC�ͽ��_��a�ڋ{Z���b�N-��$� ����͑�`����G�K|��g�.*�G�X���AL��9J��mg����X?9��bSZ܌#�&LN��xP�N����c��������;�G�֞D���n �RF��%��|�.��	��v�PD`�H��rέ�x�ڻ����A�<��=������P�~�եC��k�<�4�'R	�7��"�0y~�:�9OKâ�ʊ�1�a�z�A�(�yxf! 7�z�A.��0B
���"0��C�����*��!�q��fX�ݙKa��V{