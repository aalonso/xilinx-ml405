XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���cx�T���b��S�!��e�`��&>�q�e�_��b��h�&�f���WS��F�|�OV�ks?�n K0&Z���
g��hdL:��O"W� mM%"+4�<T���b˝�X%�Y�"�,ն�j�c�=Vβ�����=X[����1�8g�tҶ8>��0TJ��O����)�﫧�J�y����/)��x��Qڴ�Vd���H��Qh>N_�c�@%�w[=�H�
�?��q��=߫�`;8���԰᜽��5���a��;
�"��V����7t�0����o��r��lF�w����R�m��IG�3���{`�_�Y�ݜ:�]�v�öR&1�K��%�
�
ߎ�lR�$$�t%�U�~�s$��jn������j,)+�L.nw�ZK�dqҰ2�5O�v�:>��6vd�G%j�+h��"���K(c�*�VLxLC�����R�^��'(B�Nw�ȫXw���Q��L�]y��g#�tߥgJ�&�뵄lK<(��b7����85A�D�g�ȍd��Rl�~ �;�I���.����m޴IH(i�������\v�~\	���2������
�}A݊5)�g0G
���]g�;+Ȓ�{���	��y�	ۮ�/�DX}��zqh�h1'_�No���O�x��{Ղ�t�<&�M�� ��l�FSL�z��5�(K��F�6�x�U��ɳhC�Uav�o�a�n�T]�?Ə!�}��#��p*y��D~F�[�����ߗ���*��9��j�i$���_�XlxVHYEB    3292     b80� �TD�u�1<�>�'�":o��<����P��	�����$w� �j�/G�9ބ���$.8_@���J8u��L�=ۃ/���+�����B���n���g���i�LC�g �#�z�/��]����F��ӓI!KS�VX�a����}���ʛ0��L5He6����d��d�����s���Q�K�o�Iw!�nb�u
^�Sh�t|�=#Si�۶�W�����`GO��\��i+�%|�'i�x�Qq��hV��E��6"�N&q(��Z��9?�l
Xx'
�����O�v����H���Ұzz��G<N�$�ϴ�+�l�6̪����V�v5����п���WG��8I47�z=b�ж}�$2
�p��}:�~6D=��h*����P�|â"�=�D����ϫ��\Ř�d)�`���"~铎D�D��sJyY�|�c���w|�f�-��9DjL�I����g��"��3b�跖�߄���}���\B���W�c�G��o�x���~0�������Wؖ(M�K�iԅ���ĺ�;��7�e�#\�)D�$ęN�B�^��N�m��M�k0�/��m����T%�Œ7OHd����*g+��c��\���`?Lŝ�zi��{K\�,`L��§�~]�Ag_q�t�]}�� 
#��fLt��"�j�ތ�@ó��jko�ڲё���l���EX$���qS�(ր��2� ��_����;!���3�t���B�:�^�Nɶ��P�n��-Ԛ�脓�T�>�i����YZ7�٘����n�"���rd��;�\�[ɍ$��Ƅ��U���p)�.��)��s�� �.ߴ塲[���i����]0cD�IX.ά���y���g5N&�v�����6,;���,�U5f�eW�.֑O�J0�į�+��j�:B2��2���d�@oU�J��������WO0�}I�z^0�By~>\ߛ�O񰨡|��S�To�޶��>�JE�MEy�:f���:pB�6S$�!�w�;`��[͚�����'�d��d	���XQ����h���J�z[�u*`��l�oЯ��l-w��cc_kɰ}���}�]G�Ƭn1����5χ���5�����V �d 8v�s�8c�b�Z�"ԟ��i���,�f{�PII���b[C_0�+�<W�y�t�"�/�<�~�=(�cY��� 0
.!h���nc�|7)~ɱC~����f�6�(B�.��"2"K��J�	�\�%�ݿ�"�Y��t�z;Z1�>2�Q\������L�񶎔O�RpB͇�]7Q��5�~��V4ɮ��'�l"I�[��(�	��5g����5��Sj����a"��?$�6��7�7�P���vT�k��Qnu#��(���T~�V�o����u�'�ͨ.�.�=�P��E��h�����f-�
+�8^l7(R��2a3C���nK��GX��2�+���s!�F'�h�zL���l��S���R�	@܈��5��!|�0�+�]���~Ɲ\���Y�y7�ԧs��ס)����\8@��� �,��)��s��b���Ga�D�.1j��[{�q̄&��N�Vw�ᗅtv �(җYN�;[����S�1?�y�Gs8�����KABBi��e�!_;X����@pHM���-#ڙ	e��Jǐk��y��~�gԜu���9���LB*��bT�t�fލB.W�u�i�FuhK(�Dq	K�����϶�R8�$�����(:�Zw(;�����ɞ��A����N'پ!�^釸 BAs����ڊU50�X�*�\�-@�ꚨ.'������xs��{�ϖ[��L�Z�r��RD�K����u����|�|�m�T9���%!�	�n�C�_]��OW�?��5�P;+�����뜛v�A�Y�1�h��}�����A�-o5
�J8�s�j��g���S�^�<H6!1�@�Hfdu��L
հ�`k�yN�%Iw?�9���+�yd&mx�Q�N��{X�s{���^3��{�ڪ�Ƌ�4_���	4N���a�u��	pҹ����Sf�A��K��W���.z(�H�B��ܑ��p�����܊5�?p��N�kQA���ud�"����8Ef�j���Bِn^l�s�5��O֡H�*m�}.3���_+�r*+�C���v�r�@ >��Gs���
��՘:�9�ZM��w��a<�s�?������HN'l�^U�3�5/�3�G���K�.7�e��X�s�5ν`���/�h���L�7G0)	m��m�&��	^n�@�J917���Y<���2��ê'h@n|q�� G��� +�7�.����Oc���|�N�웃Q����;�E�N���=��d�uXkoYJ�T0ci�Ǡ�bA���"¹vo���,��u8��F�@8җL�뚁�)��+uN��
H�[,��|c~^d��m�+�.�y�v�"d��*Ԉ�O!���;P�s$P���F �lF��R����a�-�*y��L|�a'�J��d���ABKZ�A��z���e]����� ��P��X��5@�|�;����\a%�pF-�,8�H/�ob52�����}�\X���I����I�٣�B�BS0�`)nz�����*�UѥS���dR	�$�Z�]����.rS��vþE��N  .XR��CP�#�r�iY��A*t���."X�ͱy�Z ��#�Hv�[�Z��S������ZG��Z4r�m��+�R���@�U~]d)��@j�+����8 �9o��ν�b%�H\ r�C��:�w��z�k�H��C��F�9զ;�^�t��}��GS�o��C!{nP�H/N���I��پ��uN�#�R��u�N���5,U���p����LY�!�X�#����yO�ͭG