XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	��8A�����KҨو
ĉ�In���I�D5���=	��e��n�Y�aq+v��	����PԌ��?b��\_�n`�ᬢ%@cy�e��e{�<S�h��Vc��fo���̴�4Fi��N
r�Ƶ�m��'�rg��vQ۔?�h��{�AI 5�3��S�#1+r��)@���&=�+����(V"��q�����\[�V�S��o�S`-�'�@UO���������4�4��,�8�{�Q�� X�E)�{[v�!ƪ*�	�bzRwJ~&�����	�;�m�e��)ᙪ!���$�s�5����	���h��uW� yp��C�Ry�Jͺ��ON�'r
������_d������/���H�w����A�8E[2�?:���V����!�@�{�ф?	V?!�$n^OH����R���:�Nѽ���ͧ��C�9��Q]���#R�M;$��U���Y�*����Z�6�2`<�s���YP�m0��q�Kw<;�����������]��+té��4�����V�,�t];5�3��/�J,�*�]���F-�"�!*���fF��k����y����Ai����~��)A_93�Aͷ���B������L<���h��<c8X&��Ģ��� a+!�w�w續E#�����R+Zۀs�k!� ��k�.Ӗ��.���>�(�투|<͹9��Ѩ��������i����C����٣	�=oqWEM(9P���Pc�:6�Ep�Ϭ"�Ԩom�o�&mǣmB�H��XlxVHYEB    523b    11304c�W�b�>9�����M����";��" n���ԧ� �M)�|�M�lv�b|7��w	Â,��ٖ�A��v2�hS����*��Z�k�{(rz�0�.O����R��D?�`����d��-]�6w�T�J(E�P�F�-�̾�2���O�����][q���"g�}�*J��i�FXk鐪8XWDzɉ���l0V����9�c�%�VgmyH�嫂tO\o���ܑ"��+H}�L��^&U�^�C���D[����GD�;�4�[��P�����hK��y&�r1gQ�^T[WXҩ����n�\gMMŃ�R�-Z�o���|��7�	\k����Nvd���x�.����Z`*����S�x�������c:�G�Ð(������-�Nd]d��	_��@0/e.�3*;2�a'��dm�~jv�d�҂�_�V��S��M�ɵ��(��Ԧ�2*JB��U:��l��3H��A�_S�msn-pC���'+�CQ�m�.�/Ƒ�����>�,��یp�L��{��k�"��p�������Oa^��e$�X�
Ż��8�8��OhE�;�`G�!�ux��J`;�{�>boI?���n���z��a������.T}�DG�״��D��b�[A�y��݃l|���!ҳ�3��)�pe�h �gS�[��%��99�\�;}�A=��/��.��==qp�P">e�	9�D�:�M�mUOL긁��[��
��p�~U��-���wH�H�̂[�)duj�kgw8*Jrω�/(T� �3a�]"o�^?u a��G��R�{�<��?p[�,LhqV��&�22��QY�
Ȏ��~�a[�C��x�;ȸ��^.a�=L�@�I��KtɋG�2Agd�?��J)���o��(U@o/Ȑ�^'u��L���y���|篹DU��.P�3ٸj��
�s彈���ɹ���e
��D��NoZ���p��KWxh!��'͠Qm��ٟ` X��<�]�ߍ��,��������4z�S���F�WW��P�6�C7�7SVA�[��I�Hz̎�/����8����(?��:�mB���Ҿm������; ��}��2�zo�I��Ү��4�_�q�q��/��/'Azgv����g���_V�O6+7+����h�i�In�9�L5��sJ1��������>�m;��ҊUX[�P�
�i���2�B��sbY�&7�$�h�{���J�\���̌���F
�_b���O��g�:�
���_��9$#r�u��:�f� ��d�M{���F^Ȅa���/��ҎV�(��r�
`�@�ؼ����Nd��(�ɍw�H{3R����v�T�7��:.���cg.�ϴ�?��[�p��?�uF�V�Y�)=u8q1��b��iI�ZG$"�"̾Lxo?�F{(g����)��H02G�[!8�3��z[ �Y�I��G�pW	�U��.�_`�]��Ԝ3}"�>l^ ���N*ՖB����*���ػ�D࡛���sQ4�X�ݥʏb�:8��S���.��d�M��v�#�+����������Y�2����Y���l*�f��"+�tGe��T������7(�!�1�T��&�����F��`�
1���{��޺ �O�Ɍ�`��K<V��R�yO,���=�l:�R���*0�n�=lh�$�c���g�*ŉRTi g�|���sV�e	�L[<�����zG@�C���DN�U=$�ک|f'z�؋��,vX��k٭�O����'�)N��(�{�qHgvA8�{���0���A� �:~�p+Ë4jf��#PjY�2�W8�����6�z->;:Z'�E�s�@��+O�2�� �6���K��霷}+B#�Ԗ����jEs �l��E:�*����[��h�YB�M�h<w��y3�?
(�6�ĕhXb�5"b��Õ��ڹ}�(�x9�X�'\�3� �>����/|1�E��B��ǃ�9�Ҡ�^܏�/.ϲ\a��v=�Yd�ɘ�#2NME14Z��d��s��?/���%V�6��)����v
���1�74L��C&� �Ӯ���d0B�S�j��Nt %��q9�_�w ���UR*��鶛�\a�:x-����X���2��L����L���r;��mEN��7�3�6V��C(����h1�(�m���'�r��S�_� ~4n���R����r���A�T������k��S8di`L�=�?7�@�x�8�d����W��J�*Ҙ��Yo�x�����܎��6�p"�%��T��B���ɳ�?t,PQix�g������l�Ɗ�93�L��>qbr�؝x�G��3���<������qҖt�
!��Ovd�G�-�/�B��6�<�sWs_4H��m{�{>c5�D%�LM}����W������$��Q~��tb%4@Wd�lf?/���$����Zw�>s��<�	o}�@��C�Q�]G;)����9����@Ę�u
�G
r�˝�%6>`>�ؕ˃B&O��6]XW�F?v���[˝���̀������0/+L�ܻ^���>&ǡ[�ɸ���mr��D�i����26�lo��B��/)�����u%s|������%)�㻺W�jG���Ħ��!v���w���K��[�>�z�!�]6ܟsݣF|�y���|YU(W�b�x�脐��1�ʪ��ŧb���|���:�s]��)��E5Ϡnkl�����\��>!T�Z�M����i��0��m�E܄���⺙|NX�Au?����ά�*w&z|
������T
#�~[�HL}cykل�uǭ��8N#=M��9�V�B�,��e��ӊ�\ "\0�Ћ��1��" (dU���\��ʱ�XMF ��wx��s�z[�_��9����*��ʧ�1�=���U�pռo�W��zDp�b��5dx����O�b�E�k�������K�C����]]�9�m��oN`8(Ñ����?b���7g��H��r�ۮ.����� و�</O��]�^!c�^悙pʵU���+�}�J��X�ѫZ�v�st�:�5�us������.�Cwe�F�y$@
{�Em�ޅ@9�!��%��ٵ��SE+��"iIP�OQS�����%0}���fnl�ǅO_�덑�*(쳂
���AF� ���wZZ6�.`J�D�R}iL>=��g��%!ΉwS=�����R��,uц�9%�K	=�F�DTi���5����(�p��*��"�}�{v8�_]"��3�ќē�*�����p��y:)q��g�ud3w�X���g~�� ��P!���R��L�-`�4�3)s�sᜐ1O�v��>Sv���bu5��M���c��68�=qW}?ڀ�s�X^��F�2y(Lxx�I�Y�b�Pִ��r���O[��t}�Q'�l?�nӛP>iS�P��Q����u*a3��|c���d,�Ks�o_��)|��CZ�~u^��/2��C����<گ����!�|�����gLɆ�bX�k��ͽM%ɔZ�����bo�I��f�� ��,Ǝ�z�,)�8%1F,��G�*��6y锆���&��)k���!q�u���}|�#[���퀅�I�x�`�w�y>yT�J��)�p	�ߔY�=��f�p;�l�����Ŀ%�z�R��عG��p�o�����v� ��y=�]�-�(�:m6Z�׌��C��_�mNyb�+����|`ಔ��8�#��,�-Ƕ�[�ĸ��&�p-��5b,ݓ����w�M����\�����Ǹ�`̏��uE�nZ��+��M�k*ZA{�q�+�F&di~X��HdN�r��	�K�"��u�Ø,MPz��q��u�w��*�� -H*��|���n]�I���ȡv��j���By��ʊ\��Fc�P�=̇c�<��_��L�ﰪ����QX�h�d��\uL��9��&�����b�\�詜V�78Hãİ�Qi���TAo���h����5�x*wDrqzo�f��]�3�'�,Ԏ�ӛ3�d���#I���=����>rs";ģz��n}Wm�}�P��1ſ�^�H��;��.`���<��S��{�E���t+Q�3���]�y����	��/w�����XT0tq��=kL�&�A�����'j���ȟ�m�
�v���K���L֨�"8`
���9��_����:��ܯ��iy��� 	mFMVț\�ޞ�P7#fj,�b���b�}�3�����2����=�������_ɰ��"�.�tm�>HP��� DN�؜�9B���à]���/�0)�AL6��?黶�