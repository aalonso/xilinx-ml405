XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���H�pq�􇍓de,R���C�2��%���H�	C b�{8��=�4f��R���tO+����������m��]es��|Ih�������Xf�MO��;��⢨д2*xp�:0A�O��O�Q�f�/]@��=��XU_�q�k-�z9�4jy�3��W��rݘ�C�+֟%���S�+�T��\��T��{ζ��3_:9w�h6W~ž��C�2�m�J��$��ߚ�u��������,��s�J�م�G�5����O��_'���Ubʹ��/��n[N�4���Yk(��csk ��8����X��9 ��3��5��wӝ�:&�I��0(� ��t���mx={Ǥ�Bu�MI|�/��{ޗ�n���F�+#����u(����y�
ׇ��}�7���1:B�M��j�#�C�4��q'mHO�����qp=��l�%���M)��/Y��t��!~��%+��H�ҩ�c'������zvF���S��鸏�t#h�RF -�>��|�����6n��s���jTЛ2����n�(H)�w�Ѷ:L��樺���ȼ;����I�: ��B.�U��_b� O� �xd.?$�F�/���@�YSG"a�S���@+9��������F�����L��m��*0��S~���A3]�og1����j/7d��L��<�sa��%'��Q��� ��4�r��X���G>��A���@o@����{d���΋�L���9[%PTf����uC �R��X�XlxVHYEB    4071     db0��h#���By$���ap�4"&�
P�(�N${���� ��	Y�`��lҜS"w������!��N8�LB�hI�Q��j�U:~j7!�V�vV��t{Ge!�ў��q�Ƥ�0`H�Jƀ�&%���W���Hx�Hl.ʞ.���Pg���P&��^�<WU���}�=�Vj�ƪ�,�Tk�[����nZ"GGzoX���~E�.�C��de;�$��]��,e�Z��Q6R^Q�.?��G)�Cc��r�,���$*BW���]�m�!�W����-'hwK	���<s`��+'M��sܛ��%�$�v��������� ��7�K�,W�Ny��E���	O���/��U^{�J�=_�y��Tur<���@;�k
�$�+�V�l�֊P֮2��f��/f��Z�C��T����%�7��ڧ+|�\6^j�è.`₳@z���=�~���/,SD�tv��Hy��Е�\-6!fb[�����RV�"�dRKA�� �����4j���������J�F"63-5�R$����TŘ�3ZL{���X/�"n�R����)�.fq�z�[w��^�O=�!�$+ζUFމ.�=4�<Û�qV>N-y�J���}��A��6�("�4P	N��P]5+�Žj�|
��ij����!�C3�"�`�x gkؤnc�Z$Uxf==�W�6���C-��i�����{�Mz���c-�k�/��9;9�g�	C�����N&Ej��e��]�ڌ^�/�#^.p�D>���=�I��5�!J(���� &S�n]���"��qO�	��X����(���L{Iw����,�"a>�d����1=���Q�J�/����*�<�*��g��9��G�|�'r���y��DϷ�R����!��6�ܬ�4I�ؘ'���1��zQ���ևiv���}V���f��:Bhd�q�Ts�[�^��p���ࡈ�������&��P�G��&^��Ё;i|aFJ���Bx��ɱ+N6,XD�#(��]G�ip2)�<_%4�)��������}��]:Y&���!}����e!�n��H��$�����8?�$�v�q�]W'��O>�H���n�Kak.�����w_7��MU
�J��a�RX�l�F�H��ȮǶ�4i�}�ʣc����ݭt}8$��(<|U}I�M�D'�T��F��~S3�C ���i��v@���d�� ��]����o�}��i����F(E��u�S�������I�T�ͱ�xoӘWs ��Y^�[J���$t���h���	U̗���L�+?G�Wa宧�B��^YCn�0G�Y�ن�#|}��ŵ�j�0f�&�$_X�"!e��qCC�+ex�N�T�)�s�Wt�T�a�s>P
J%"�Mb��^��t��.Jl�s�r��U��m�^����@2e>8��t�nz��EԜ<}weL٤�y�E����v��a���"��o~Ø^݄����>�9p��)�L��<�|ԺcTg=WJ���L�`�7;K�F6�#�� ���2�RSf�T_�W$�2H�(}��6����zYET�+kL�'�a�_Ae���?_!o`q�F�8�Py����ABh�`����ISAɔ�.0�+��<S����ip�"#!�Λ.;��,��L��rH�00r�(����N��BM�̜�d/�ID���"�\��;@'WWv���TZy[ۉ�w����G~���TO(�b:ɺ��a9K�a�a�v�ﳂ�^�k���z.v�����JŏQH˽�$��J���)�*���y?�
c8A�O�t6R6�&��.Ź��=���b�tN���+�;�}w.�:��M4e60���L�"�U��TB�1Q*�tN���͌�s���� ����fbOd�_�r~�E�'%��������5�|�ߎ�S&&��fW�1"�����U4����H��	V��тS�4��Ij벫�$�#O��	]�[�F'Ĳ5ǒv9&�Ne�c["��e&�?M��D�B�:,�7���tEV�VG�=��=�#?;��<:�8�����3�S� �G�4$"��L4�SuB_S2TB��F�Eg��2?q��q�߬7y`��);�y �* RŬM�:fף��ZS���,ͪ�#�9�DW7;�]����k��x���� ༡���	xB��=ujn�]2�A$�2G�&-�\* �4�t����X$}`|� H��M��>ކ����V��v���]+�,{R)��yeg�|?Q�p�ҏQ�y�a�3>x?5�V�@K�=�K}���2�-�����@Z����9���R��W��-b[� `+��dD����)4��U��i�R��T������ɣO�uN�⑥�,!F�� ��+ۑ�mlA�a����v��
X�Ib�8$i�`�UܲV�M>��Ւ��A�0���d�X���R�M��u}��F=����E�3��~^�+RH��	wT�A"핥�_��ߞ�&B��'�5W���oto|Wh%X�oC&�3�̊�p>���1�5�S������A{����PŪ	O��?�J�'��W��Q���Uu�qB�d�2;3��$�2	Ik�]V�j���эV|+d��B�2��{��	�g�ߡ�*��,�##	�����@_t2mHi�_�nL	�o��OF�V�cl���*������5WS6KV�)G嗨��<QH���w��ۢ�x�*�[��ԾU�O��jbVEX������!ؾ'�⫾�ۿ�r�����-�|E��S���)8��%�	�Co�=M��fN )y�끊����t<qk��V#�7��,&2^��L�w��l06Њ�V�5��O�go�y="��q�F>�x��U��%5��i�F������pm��t��S,��f��xP�5����!��C��?�F
Q�J8��z�7�y�z�k�ڢ����}%Ϯeʮ�aE�vQ�v���|2U��M�_��-�ђ��|J�#l]�/�f�kx�Qe\%C�N��E-���A��&a0��]l܅�+6�K�H���md'�q���aN�-�/8�ǩK�iҲ �I
�O�%)b.9=�A�zsq����hc@�h�b���L�q��Sx2��M�xV�7! �&OѾ#گռ^	=�8��q�F[�m�
���ee��.�@H
o. �����2�߮g|t�A�U��EP�a�"�$[�p�K�? o��q演����R3�N+�v,FQB�&�_¿�*��k��̨�߀���H�_Q~�M�j:df���������R��}y�U^1�.���3�V>O�@�#X	</ȡ�gߥà�U�R����`��5D
TY!�Dk�� %]"�.n�[���*�q�2�M1�E����RFޙ��V�K��P�&û���8YV �Q��m��g����L�����1Bc�0`i�+�ȵv\��}N�)q�c3�����[7�IE�����:���y�