XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?v�G�Qp,�����u��ӟ��� ��n���Pr5��N+.{� z���g֤�cay!�$�=� [&\+�#9F ů�H�駵�]���Y��zU��4K�
�|�G
��ˎ�G_�>�QZk�8u�d��g�����R�.&�����u?�:L�uj��k�#��V*>��hr<�R�&TB��Q��ԯ �R0�M������(bn���}�'it�Z��t�")Ja���ޘ�uGHVS���|���8Ơ�	&ݛ���;�)0�0�ol&��6VN�� �Rs�li�&K�|Cp�h�.����هi�<�rGU<ҝ��j�w����k�����&�:�6(,r�d
O�٤3������l}�	gހ�n�Q�������*Z�q�T�ȟ�XG��#��%K��-�5UӰl\�;��� ���>��n�* &������u�P�MQ��p$�H�>W@�b��B����]�D��b�G?�fi"��ऊsg\�Y�һ��WZ�5n3j�cH\��z"6��^BTL�9�ט�U�������2ſ;���W�����9_GJ�C;)T�����e�»�0���ҩ�K�����#�H��yg�L�ᝄ6I/T�����?�<��:��.���W;��צ4P�����tADt��&v�h�����)E�yI�|I�{z+���Koa��Æ�	20%˴P���M_��1�Au��)��&�g���XkI�9����"�k����_�XlxVHYEB    1231     7c0�J*'�o�P#ޡ��OtFQ��z?H�lM4r�'�3t�\��0]��q�Y��i��E��Q� �J3WBu/� l�uѝ��ù��U�y� ��B\q�i����Q;�?����F!-҃DA�o�v�W��{FU������+���xx�'G�F�t���̢5��jC;G��s�Zb?[���O�51�j����U�M��yN�S�!�Y�k�V�� �vm��6Y���D�^QN�@�V�圠UK5��ɩ%u�R�'�-�a3��W���>��(] ������~�H��}��L$�\��y����j�����C �*�}��V9���2���o��W�X��5jl�.Q��s��īp?s��;<,߬��۬=���eg'R?Ѐ7�8i����*�I��u��z�zT�ѯ�qo$�����bZ����(� P
���H@�{�A[�'~-�(C��>��RE{6Z#�6�u�15�,��M�ZFY+��=>�_�_.�v1��~�2�Ӯv墬�ga�#�s1�v�%L����~F��b����8�����m{�î��T�\��?���:���[�x��r\,M$Aw=�:���j6���J�{V�L�j���B�,��"�4��E?��0{�&��{v��q��K ���;��앭��"RN=������B��&�o/�+�
�\q^w���Zn���軂X5�	�}�9dن#C�f6�LW4��L!�c/��l;k����v-@ժ��ޔQZ�;�t��}�g	lDOs���S^eSg+�S�-X�_(Ęt�N��W�l2�	7���nu�;?@;+��?�&h

F�9��z�����;���t境���h�L�8=�j�{�4�l�N���O���@"��5`at�G'�)�v��k}Uõ
L.���zaɬx�:��:�P�;�<ؠ����#�|�ȘGբ���m�p\g�+���U-��B�����/0OC�^[�������6h�	.���w�%�H� �1��F�<h���ֵudN������*�x[��r��D)�R��n	�Z+ч�l>E�|U�H���IQn��(>z����裛ƭ�`@�Bd��I<�X%4H=�%_� c��������;l R�B-2f���IZ#�.����7�DA�H����O��i Ir��ͭ��������[�� l۪�nt#��*��Z���4ɂ�R�:�l:��	L�1r�K2�)x;{�-��I��m�b���[�44Y<h�?������nL�צ�(��{�nz&3R<i\@��,���#��A��(2��(��|C���FxԾ��m ȓly3�}8��_ݻdI�L�]/䡖yc`H~�E$X�O����ȫ��@^�]�N�X�E��Q�a��)5�K��G=�h�wu�ѥ��H�Q=�1l~��@�5����䢞ĜYxDYf ��`R����t,T
��c�*�r)1�-[��WX6�R�پ��P��Kɼ�W�L���̧���2�t�f1m���z����!�~����\8�+��P^h����jf������JYU��
�	· �y��$��:�˓D ��[�AC��\N�����*�j�ҢcyQ������&��ְ�p���j������å�hT�d6��3�$\ەJ��<xH�2x}Oн����]!`j�a��f�63����+�lٗd]�c2����h�fG&�gtHƄ�0t�T�ʩw#�&�v���$sJ�pȰ(�'��uM�{�vZD@�򵜷ot�}]@bVm��%�ZW/�4?8�c\b��#�L� ��W�`���(���P!i��g �C[)�/|��Ԝ�]n>s��*���:��e��\N['�B�?�3��H9`ܚSz~��3��Y�㓂N1�;��Y����?�$�)��yF�����S��6o�����%V����l��B��p�1L(��y��#���5�