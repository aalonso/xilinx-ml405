XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���m�Ѹ��B����*�^!�6�f�D�*�jS��7=]=W*���%�%��CWm_�.s��0r��ǮrTK�*��!U���e8R���`#�8�>\Ǟ�`��7b����ϥ(P/��ҍ��ԘB^f��}7�c2Z�W�{�U�hn��m_�Gg�3ux��5n*�'�B��z[� n����c{�
����;|0|��$�˔�%:�1��[�^��N��#�Vw�u�	Đ_B�{}L}�ڈ!�n�)n&���p����Q��N���]t �b��X
dIĭ��9��DԂԌl� �uHwٗ�3Ѓ3W����~�WnBy�~���"��`5� �3���1�$�j��Z�x`�#�������V��TTt����{	�+���$�Ӥq�t�)�g�_��TsC"-� ��@�u���"j&r��gFݖ��ʇ"S��,8���<�_��Ǖb?HҩB�ǰeǚ�c�.ͼ��vL\��v��ٵ�l)��YSq�I���/�Ԭ�;��]��-T�mg�,�h��e�a]��	I�2Q6�i�b���_�"'��aN�ASG*���h��w�Z^�bw��2�3�D�qGy`9lZ��D8.[�}\���*���=��E>|)�����t1�O.8�$[�~M�(�>R�P+�)��,��&�Ȣ�bl��Y�6vR���H^�t/�+�{��"~*H�:a)x�Ȓ��4+.��hn�Ks��m�;cD��!�-"7v�T�� @�XlxVHYEB    18fe     880����t_h���S����VDr���B@Y�/3T�R4�9��q�xrRf�C�K��=		7jww���P,j�4�F����oe�1������@�Ou��S;�g����]���
��y2Tl���ҬWөi=�[�gL�����`�1���e*�у�����ͮ8���2\�rz=	��[a���F��c��o�0X��Y>u_����(��q�peu�2V"Mb��S�'�og&������A=ӹ����0���al�nj��t�UGf/3l��
e���P'�9� ��~���_z<Z�N�|N��`�mojkM�V�q <>���0�y3D0��?r�3�8઱=86��1�N�פ���-��	�����~�<���o��̦��L[}k�oy2��l�<A��������9jϜV��X7o�j��4Kx���8�/4񗃟�|�,� ;�!'f��L����!���
|���8��_����ol���	�l�h�ө��y��)��l��̧�����zM�'♖��3� U&���_�pE9;u�mq��i̈́%q�v�*���fQ#y���Sb�7y��[��s�����4��I7��KH'�s�9MA�q,�>��!߯�l�i&�Ae�Q/�-��A�'-��?Dΐ�ɕ0�7��� #\]��5ָ�@M��Rh�M����e5��x;��J�&��B�ߛv��@]hX��F[��4����G�L��7�Bd7����Vi9��3u=q�0�l2Y̐pBע6���|�Z���(yU�_v�~�.�F��T�h��n�Uɻ���V�s��C ����	�-_��>m,�T,7������G��n��l=r���rP!w��J�Q����4K-�M!|��5�q�{�H�W���x�7w���^��J#$$������`��E�@ؑE�H\'��z;�/��~4��H��%��ldEk��7�Jb��:���E�����2I3�8D�בq�m��4A�.����V�;�U���_D���x1������u���[���8j���
tpĻ�iE��A�ww���,ڵ�;�7���D�[%	�d�ݵ{�(�ܸ�}��^��ܔ���+�ýV�ّ�kT��jM!��I�+�-�{U")c�S/)�{����J�9�Q�o�l%֑l��p�G��%2������8iõ�@�h��U����JC
��y�
�[��׶+ln�� jy����ӭ m��՛���
�@#\19��gs��t�'C*�6�+��]��F'��^��j�>�˦w| ��vX~��]|rn%N�A�ͣ���"��.X[:Ը�t\�d�P� �"|猩z��o=����!��q�`�/�bqm�8�v)�X�棌���ae�F%H����m$��5����^7�/�Cƹ6��r6�#���-H�0��#�^�P�k���!�5%dw�����8E��_�mmq?�&��2,T��fN�OJ�	^�Y���y�*c{�cxqdXö!�1��g�kIR.F���o۲"�<�n++~�|`Bl��=��Eaz�OZO��qH�G�L��3�Pu{���w+ۇ_�s���(���0b�T��V2&U�,�WE��}ė�,���T]&K�I!g����9|R�{U�;}	�m�>:b	��������7T6!�Gc�5���H9ð�Cw��u�Pr3��s����?�K���a��O��>�"���F5v�� ��*���QmF�V�ʇ@g����ޠ�Eѷ$,	T&��w �J,X{<$}'��`���9��4�`��J������>E�{>�lQN+�����SN�j=�$Ak3�?�o�]$�&��U�cS�C�.;���T��������q0F^���%I���)D��ڵ�Us�i��ׇYI��)x˧!����䶒��I,����=�[�^��'ҿܦ�D�^�n��L�&�jK�;--�?�f���҂B|��E���H�J07��m�ԷRu�����l���Y�u�̌ l��(p�h�'��+P�;Y3I"ѽ=��:Npm���*���87[>[��ĺ@�/�$c.K>}"M��2�*��Nq)�͑�[>Nn���2!��rc�{�HB6���S�m4JU䘹�"���xP%��?��n�#�-���bG�?��U&�|�