XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��>�Z��:_��}�)H,�yX����N��njMɛ��4��^m�<rod�����Yۥ����@�LQ%:{߇r�ۢ���WQ�f�ֿIf��]ނs��?�'��5pvϟ='~ ��C�٪O��C��:���m�E3�'P�.�Es!�� "4�G<�4::�A���A���$�e��� #�O�:��/������?3����D�aZㄭO�M�ND|X�K�92e�������wa���XB=H��m���<�yz���V��끠>ܙ'S�<��ٵ"�?W��0/о���B�W-�e(����Ƞ;�H�.���Z�Ԏ���$��T�E��}!��.=�#�)�[����L�9
x�(y��5$�2&�ӎ@/�#���(L��0��V ��a�C$��EP���T�eӯ�Ǘ���'ZIW�E����+\�Lݫ�?��g�)�,[�%,l�pj���l�۟G��󘰷R��Xa]�n9����Iu�� �������H��`(���Yw5+�(o����p\�ɘ�+zm��vF5g^�$l4�'�"��0u���G=�c��W�4��R+q�q����"f�o�����=��g���p����͐K��$mg����Av�×��wȴw�'Rq��r��t{3�	V�6��%�����ﺢ�P��{�Ա59Hi\�Ӕ
3���DX^����j7^�B��ρ����>��}Ӌ�w��˰~w	�0���2�G5l��w80��t����8�"�y�RQ�m�
^mw�XlxVHYEB    5fd1    1710b:% 1�=i�b���d�gd�Z�|��|?י�{S45x{'�D���
^�����f8�Є�H%[�b���Nǥ�N�LsԔ�������s@/'*w�W����w�U���C�����u���4�6m��9�1�G)O�;?Q��ч�&�ʕp���� I����+M�'��~�������~�t���"�G�|��?��4��]�f����Y����K8���!���琒N�'�_"@��5��fo�'Y!ii5BZ�w��C�������rDM$���Ɂ�.��j�@N�OvŠ�A� ��3IS:B���/��%"]
��8����-
����#,�Q��D�RyMT�-�9���ed#�*������#��F���������!ӜεCT����>W0b�X��Rn~�+b�Y��urЂ���I���5Ɋ���G�3;�e�,��Y�zܙ�r>�C5�}\6}rq��l��1׋����̑|���yF��'�jd���jAa�r^=肇�w�ھ�Ġɛn�2���9T[$�*���&�^��A^K`2Tz���>�[T��c�s�/�&8Y���	�R�4��#��
��Rӗ�b�Q���V'�y�_џH�2uY腲�:����1Ɏ���V-�<{�2BwQ@*Q�/�o�g�܃đ�_�~=|�""�%2�k9�m�����`�ed�Њ��4���R��-¿I��.��Z���'��Fl_�{@��_/³3S�<�sЃ�w�p�X�� S_�JwQR�@VJQ'���H!o���e�{��� �q�4�k��҈��E�Nu�};�}��s���_ ����\���u"�:��޳���8O��ED�S�$�s�R՟�¥h��t^yl��<v�7ϩ���r�J��x5��"`w"�f��,#�k�?R]7���彠�%:"]�w.�	��
�
 V��_�J���A������ݑ���pHs�W!��Q+1	��Z~�'Q���d�t�0��U�J��3;)/���z�����u6P��-p�� X�(�#��")+_�;jlb�YUspP�Pr�O37�&hw�xY��̡̈��u0�h�b�r�]C V��G���k/=�GB�8,9�J�O-�������81����V���d��;r��iG�;SG�H�Y"��Ĉ~�&.��N_�8!��a�2g���]ʔZ�JQ���8y·�X�׍�M_�Pz���c�|Q��M�6HZ���'�WA���̹�G-ݳ�)�������b��w��eZ˯U�mz�S`�q��#�I��/�1G��8b:)��2�3�l��n��K�9��#�j��R�����te�'�.� ����R�7f\;J�2%X2!:j�Tq�KwSi��59HE�!}Vj��
D�����և;"���m���J� :b4�vR,g��P����d��w�i������2�'�O���� \��3�23�c�p�
*��;v&�i%>M���ZWP�io�ថ��l<�XXR�o�3�ķd
��7�m�VlNj�U���NF�$�#�ꉆ2���>6��
���������B�9� $�
�726�];z�S1 �S{4���d�%���i����y�C�Q0�n��k�)���
}T�6���6l%aG�GX)<���0=�x){BވS�G�v=ij����;����P{��c`�ɾ
�r�ǲ`ٸK��IU���k�� Y*ˇ�uoW������zja���C��:����r��R�k����w�m�&�����.�j^*q�=��X+�e΃A��s��{7BO[E�$%����<y�{���7ȅ�X�_�k���+^�Hx~�s��3k��)ύr4t@%&j?~ܧ�37������ �l�+��o�Ŭ��n3�4���s�&�w�<�uE�2�6��5��&s؜��Q�u'+$��2�2D~��Ft����U�p�fr��!�k�Z�[L��J�$�aN�`���z�Fl�bS��?�+=�
�V��M��|L�~�"
J���?�����S5��l�HN�����0�`��4�����23�9�I��_��>?�N���/(V�ick��Y�l�P���&J���Uw�w'�M}^a������T9���[�67���E����z���<0$F��+�7o(+��;������a��穳5|�&�X���V��1�܂xO;��K­�<�SJ�T/kܪW>�,� �.ۆ5n}�8>�	>��G���`��@Q�WR{�i�=�NČ�I��	�~TI!��Hk4צ��su `s�~9�r�L���}z�d���;i��۬����K��'���W���ejx�("�^�a� ��u/�d��:�eb܍�.���<������s_�Nۦ��T{�v�VC�Z���KQ*�3��
ѵ��_I%�1/�rd��ځ�w>A7��h�Oı����Ρ���▬�i��/���U�x���z���t��1� 6�7�}@�\8Q��8��P�ct2<���ܙ��ӑs��{�E���BS�6�Y5�H�,i�L�ܠ�x���;���yx� $u�ט��/�e�_Gc��xb��4@�-{:F�F�*�]ϝiM_KPd�L�T��o�����ۘq7�o�e�;�ɺv���'�����<:����x�3ߑA�l��]�짢ܻ�BǙUή� �"��4ʑ��J�m����a~��I��뺆
��I}�Q�B@[�!�k��q�e�j��6�A���BB������$�Ț�H$	���>�wR��5E�U]3��冋�f�9�m8����g�6Q����ژ6]V>����?��l���0$�;��}�kP#x8�O�+��V�9olD3�T+�rSc<X�;/�_�������}N[������q0���8y���f�+��D��(��L�}���X&2�b�ek_�w=��ϐ����1�|�b�9*u!��y�X���y%���ļy`�����4B=y�6��5��Ь[5����`�ޙ��зʯj!�L�k@jB%�"ѧ�EL��!�Ѫ��-(�m�M�;" �fmX��O�x�}�s��A���:�h�H��M�z��I��1���-4x���C5���
S�s��5�B���qyf7����������h6(g�������$^�f��pX!�슭2��i||D-�q�Y>;��6�,/�OEЮ�\�y�^�_|��hx�(ej�kY�s�8�y��d�^`��-!�������;�L��d ���hĉ���c�/��k6�S� ���!�}�pe9[�b�&�ސW����Q�{��a��ݤ�ʫ�iUm�.���6��cE��iU஢��m��6�t��'��n�X\ׅbo*��(���Մ2�a��Y6�Α�e�<�$�ػ�ߜ>,�=��-IU�)�-��T��p��b�c�bՅ����������أh�A��@[�m"����n�]�`�c�R�6
w���J$���y�}/��u,"���I�S�c�r}}Z8侖g8N�� l��v�@˺�� ���x�'�l���Bݏ�
�>>Y��,7�h9���ˎ���G��~023��ϾsH����ʮ�oۧ�7z'dAy����7���$��m�Hp�`^$�+��W������.@���\]�g�i��4R��m�n*���6eѦ)G\ҝi�\j�3�ia��ٱ���ℛq���>��dl~�N����%�C;]�;���H��M��U��^�e���e?��K�Р�9���Ի�x1�h���Z�%v2����wy'�k�N��󓽈)�9P����3ބ��g~i9�ko���Ma8��Sy�@W��@W��:����a�,�<��\�}���y���Q�Y5�\k�Su�R��鸯1�C��	Qt�P�&�^A� R��f�
4z%f��K����5�7�p�~�L�3�P��q�='C�1����
3{2*���ʢ,3"��1}���/3P���9��r�^����w*�J���T*���i��~9NL��=�O�i��K�����i(~D�p���(�nlx�MI�X�x����+�Tӂ��p p`����(�It	���j%u�O�Q7a����ݍ� \����Ė 7�s>��^�G��z�(
ʸ�^��W,FxE6���CC����̱њOJt�X�B��u��%L�"���l~Vh�&'50:_����b��rV&M<��'�tO�g�(�y�Lzl�go��F�+�_va^�SXĒ��8vQ�����)z�="筃�R�/�K�?܀�ǹ�'��J-��p)��98"�,`�Ŧ�"GQ����,�o9�GS��`��o��/�Q��O�hA1԰t�g����k�d���������(w�%����쏵D�}x�5��5[��?��1���	V<��}��?��_���=y���m�n�8A�J[VE���R}��8�$[��2��ɎEؗ� ����MrW�G���G4����u����e��l�u4m5!]H݃(��s͵���
�|��|	���Ь�kYQ���m,�p���|.(܅k��fK�h�d"����}}�cW��?�J�:$�R��^�t���:ŏ��~�F��*v?P4j��@���0�f��8� �O6�q<�㊷�.=yLp�Css]Q?��]9���mO��GQ���g��Ǖ�ǻ��^4E��	�	���V�=}�VS�(��;7gϚ�ٙ	p�u��~[70O���#��E���ڥ5���S!�S�6�9����&0L w�}�hy�g�����u�V}xj0�7� �"H��l!�G�T���j���I[I6�w�����]OC����ύ�{��p��x��?n%���X���V6%MOR�g,�~��ҿ����9�_�|��f��a��,|7G$��ϨRy�,qoh l��"���OW��䩉 lC���l\�$s���>��D�ŗ���S;-,��r�-���6j��:��k���3F��^h��Y�Y�ú/&'�� j:W�+�M��]Sƽ�v*�6��t
�?��|H=!H���E��Q�Ǚ1�/����V�>�#��Gݹ�G��E�5�s��Q
�����w �Ç�-�0H��jd��-m	Be6���G�ezͦ"��#�U�5�L���a�8>�ڌ�TVF�i�a����2�v
T5���$�t$�#�8~�y~�&��9��:_74#-��Q��wV����1!jp���`ߤ����ºb��aD0��DmA�d�R
2��{��υ�+�[f�S�(�!g�[��=>:u6��U��F��0h��֕���b|�V$��q��+��k��:��*$��.�����sF��'嬇̏�8ġ�#�����?�{����@��J�ᐅ��1ܯȝA*���]��g�L}��(�'���3u�����$�Ȳ`��!��l���.�X�?f�qj��s%>y��_�W�W�x�b��Ɵʻc�n*��y��o���K�1�: ���;���[e�9�JƼ���.Pũ�q'��K�8�<�����n������L�b�4.�A�?�`ku+&�V����($̑y)�P�ծ�:͑{����+r���9`�7�I���{����K�J�OÒ��������7��.���j-�����OG����H���e�_j+�\�~�D��{\*�rT���4up�M͑�_�w��k���L�HooI<{ƏOym��=#�,���'`�%6e�9�M�Q)"W�V�#���>q�י�M���?C���#�#Hg�G��J��ƥ�LY*sB����$����'�Fcv��ѵv=�������	��ğ�����-��^�?�y�