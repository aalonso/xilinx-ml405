XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b��u;�.�n��Z���Ⱥ��Ť�v�:)�p��uFG�"�?���٩Mh�^/��w+�T�sǱ��Vc�'��(�2�:_�ߛR����h	��VY�q��{�{2�f�u	1��ы���u�(>�=C7w������Mc�{q�N��U�W��������rb����<g�/g���[^��:�>���N��<Z} [̦'�F?o%�G�L�Ql���}*b.�*�8�ޡ|���Ѷz�ڬ(���-��%O�����W){5haΥ�5�H��H3����@E:?��_I�W�k2D�� ɼ�>�h��ח�6{�*�!V��V{t����>��M�La��>���RY�N���J�דv��s-��)��|�fJ�y�v����Z��ЋZ�Uoi��e�%x�봷��Q]&��!W�m����£H5�3��z��� ���j��"�n-]��ڡN��d�������YU����]jB��>��������I{����Ŧ_���@n��┐�M�i#e�:`� �����U�١�0	9���L�w}[&xV�2 7&�A��.������Ւ�g-♀�_������݆a�Ӫ�8ѻƖ�Ɛ��s>�ȍU��f5kө�u�A%h�:?���2��{�n�j���'n&6���ZI�Ӱ/�˞F-+^j�o^�@����Bb�=¼f�u^"����2�QIŅ�ނ���)Q�H#c��*^U�l�(�E+�$��S�T��?�l���O��*D��@QXlxVHYEB    d81f    26f0�M�Ry���y���;��q��׻tS��(�y��FIcG\`g��{���Q628<v$.�������d�bzQ(��[o;q����F4q37�9�	���Û��<u\h�f��,/2SEa!9���Ƒ�IC�c�ry'�ml4*�F[�Y�^��|	}���5��R���b����4T(�N����_�U���1���j�"wL@���@��{��1��M��N���E���=������d�8��8k{����_����|��8�Dd�l��?�VF;�y[��-3Fi�<�_�1���)�h5{rR	]=cz�(��k���b|�t֔R>dȀN�5��a�A!���
-'�O��G��T(e�&��!W���ϣ|�)4x��vY�q@���#e�@g�}1u 6��!�?�[�y�ˬ��v�${�h�]�bZ�n��r�$�]��kn��}�����n,�^O���*r�0n������oL�&ႴP8w��|�܆� \Kj�q��S�o�x^��jY�:�䲖��8=,��W�K�)'�3�6�������6K�}|Rc�@'��bq�	���Ҳy�YqEFٻ���#<Ʉ�ʍ|qd�JKG���ͼշp=ڭ�.�Wړ
�B�610�%V'H�Z�ᢸ~��gM���ziS�j�6y��J�w*J�a�M�+�iM4-�p@C�~��Ґ�&���ЯsX�;e�A�s��Mx�W꫄�@��^�[�������[�cb���DC�5�΄B/�i;1#~�,'�y \b��j#�̍��4�p�rY�>��7#f晳+�0!0J����@�c�q�)���������5R%A�~>9
U��g8��t�ʷ��d̢Ƹ�'��c���u�F�h� �P�gˀz���*@��CD�;�G�Έ�$1D�K�<�Y��g8M�&E�Wb/v�BU��p����z-Oh�њ�u�	��#��YH�9{��H��`�.A��^zV�҈_��'d��"P�47�Y��S��"s�0�_Ě$�)-_ŧ��	l��{�?�aW���*/����m����<��ڙov;} #���V��?كV�-�U�d��G��Ȗ��i��o��qD4@��jvx�8�`��m?��k�~�`2R�%pB�hY@�*���(N���R��$��4FI�v���	'�)#u�kG("�/{=�a�� �W��l�&�K�U ��(��B�V�(�=��#=(Q����o�Ck��ژ�K��u
����U��f:P�.�~x���D�Z��H>��#�@���,��]"�z��a��gzv�#������~���]�φ�EM(1�j(��G0�ƚo{="[Ɗ�M�h,��Ym�>/�'�:��m��� ����*��x��d1\aCrT63�@��@_r��������G7��nR�6�U���ʡ6�f��������,]dI�q��8aU��P�$T߆7Ϧ?j���#�i�Ӻ��8	�0<a�2K_��i�p.��%���\����IV��ar�CB�m�[���HYn!���y��[u�嘥kZGa�)��[z2d�=$�I\���~��Y��$K���_�����҇��\+Kx��%Jd3��>�BQ�ej��/���J18$}@�GO �|%��2IN|����MP�2	�p�f��!��fѓ�(�#]�o�F����S-��M]*VvYT��ztɦ�z�R����Qw%�}n���1�����R��[󭹲����2���3(��@�G����'���-�\�Pm;�2�`�y�Y���t/�R��H5����[�F�=(ٺ��Ӓa��9�����)v�&�]D��i)����Tt\滙!������zqP;U�t���� <���!qh(62T�.�^��U[T���=����㸆7Q�#�w�i5Ѵ�h�}�}��+T�( V j�A�����*� � ����|���
�h���4Z�g�p�}��3#C����'o# �U8���u�)�d�߸x��n/�w��!׋|Bd>�aB�E/����ٜt�� ���e&�����Wafh�!��rd�K����}Ո� P¨њ��
'?+�MO��E���Wo��|��|d֥=�m������ʤ�r�^Y��~��H	���� ?�GQ����s��K=���w �������a��	�lG��T+㮝N#��H��SC�׵�������U�-�8`i����Z�w�AW���ze�f���4+���@&|�sr����4�Xx����^����7����G�y-8
(��eDbS�ٵ�Fo:���<.�ĝ���@�ᣭe��챵�����P��n�5�|���g��Y���[�a%̢�}�᦬����aH���C^�Yך�-��%�.Ԯ!I��v�i~O�jԢ3FVQYS+����Ƭ*=�d���
�>��E�`����(d��Y�z�Z�����kU�M��yػD&x�]�E�G������}6Q
�
g���$Ś�~��C?ƚBMJg4@��@FX�z���+}����s��k\)���|�D�J�-�8�ɟ0
O��%���׌w���ݯM� zv@�ܾ.ȩFo'I"�O��M��"�T���;�'P0�)�`��@Z�P	K%=B&�؍6���P[{ߩ�""SѕFX=�Y4���se��M h�����q��M���z�U�u1�먴�Ȟ=�k��i�#V�L5Y��e�$��nE�y�S�1s�e6'7qc�E���:ğz�Ŗ����K�~r?�/<pP��Ha�N��~ⵦ]�,�UK���HA�]t�M�[D���6��Y�emG�j�uK�k9����J���{_�'�'IOg��ƭ1��.����Y�p�P/����p��u$P,��S�]�g��H�@fa�l���_��篾�9:��B,��fA�M��n.��,TE���]eN�{E���4y׼�0�R��B��$<�ބ�`��<�T�w�$z'"��EZ�jRo�W�%5�G��d��K�'�v�0�8��Kߡ�>���lD6�\�|3��DțU�|'an'����J��ew�i2���A8�x3��<'#{�k)+�O���(�m����X@M_�V�E�2� ȕ�]���,�Yae�?��jS�P��������}\�uM��c_� vEΦ3MQ��kr��(!�� S�
���.><mI8�gZ{L]��ԄG7&��J� �z�g@㳀�a�����-��� %�J4����0����eq���N+>�󻚛��	G�*��p�Zv��.�6��@������t��|o+(�y�K�4h�(��Ե���_�d5���N��+����G<Hx�L�� ���҄ΩϘ��yM�Ip��X�.Y������ځQׂ_V����<[Жm���JT�w���D�ª*U���>��+r��r���`�	đn�Zf�/���;�<\c�iD2��T{��q��=��3�Qm�B�p ��F�Dx��n3l�]M#(����(-�$ֹ�YI���p����G!��!��[Dkئ�g���X�(C^�ʲB���}��Tqq�Q	�~��O����q���iugJ�?���G�d3>�h��>�\N��/e�
�5TY�o"曧O���eFUNF\%�xq�g��x���p!阞5��e#ɂD���rK���v�� b j����	�b��[�iKa䓞��_Z@j&uo�U?�z�RS!�ۥ�5�^!���]`ʿ��t�l�@&L�fVPU�{�=(gPq��i�vM#O�0��x���/��T1���r�w�)���r���D,� �L`��Z�N������xp&�j@fľ�i�����O;��9���Y�z�T� �;Bi��C�p+u�Dc�$�H�C%��� } =� (eX��~��`S��Ҕ���FOh��Z��m��P5R
�o�#3�O@��P�%�Ow�DU���O/德��6�=�悛�I�5
�P��{���Y0,���V�\������3-ϊO���V"�s�� 7���~n8:f/t�-=��"��ł�0 �6>E�5P�H�i�)��6��r�Ȟ�S�e(E��<���-�󙰓�0���N=�n� ɯ�q�-KrWZ�	���h���zy+��=2�����X6��=�6k��r��Y�o��7�2՟	���4:Y8���E-���bz�����ڠ�G�D��I"��N��Zh�q�?[G&�aU ���7�5]W�-��?d�?�R����M�͏c9�*�;m �.���h���+�&��ЇD��zRx�MHt�Z��_�6�u�c����5KJDz��uӉ��Ͱ����k+�q,�/�p� �[�.� �4�[p����j+_W:�o~.�V`aW%	s(�d��?V1|Y�d �`x��茅i%�D~��=*���lO(T�fM)���Tp��J�О��,F	~�*��6OM*�;׊�D�"�)�zQr��~8KӱV_|ӻUY���'獜���m��e�SEh��-��A5厐�h�$�Hdw����,�E�j�D' �	q�měD�������F9<����_�Z���ԓ�������V�T,��(�K�;�>LN�l�	�>tQ:O��4)35K>��o_��<%f$�Pb�����ܫ���zh�*��σ�-<�;3���;f�s�ޘ���}�����ڧݮ�b���[�)���D�?/������Og�f$m;�����A	�{%����7�g�F��ʫˁL��+�i&����h ��Y$8��/�(-�砡��{�R����}�z��>��\r~�QM'�m�C�vς�������w8�����d��|	���/����D���?ס�u��}�_��Ux}��9J{�_�����X/�*P�O��~���~��z��ͪ�!9����߂���B�)ظ��eӿ�a�+�	�62^}��Q�`gu� Z��@�$�wNa�@pR^ '�q�Sg�PQP6��М�5� `�ǔ��W�ewJ�%,���ě�P�ЄLQ��H���\tT�ϐg�v�>Ki�+��A��l��|-�n��e�ur��<����h��{�~��:���y��L�>p)3��-`Hy��b��Zo#�����]K�5=�6�k�BQ0f* �$w�7�¦dL�m�-v�w��o �l:��#D#�{����;�:�*tvSNv�r��,�Y�G�Jg:�����d����My6S18N������HI�|Xj�H�3K�I5
�kVN�!���B�����ϙ���Vf�P��H����ʪ�$a�� u�i� ��&�b�J��[�3�t/�����m���%��z�3��Yq�##GH�<!4��i ӿ�@�/���I�q1�0��+����:���>-:�^���|kB���&��0:�ڎ�!C����E�h��^������p��_�j쵊�F�>�~�|oR�A6O�	`3V	�ۏ�9����{皌|�Wh����0���S��g�)��;������J�d�'\ ~���8�����AFX�7U@��4+M�~��[4�a��98�����'�jY�	��XP����9���==��+����ψȳ|.a���P��<�{�M�;G���p����w����#aI�il� ثH(�O��7��8!q2��^���6����K�|8���x���dG�n��.b�XIj�9��L���?�t�o)[_d���뚙���s��ܣtw._4�)�)��~���)�Y��[S Oi3�ZlU�:�A�zxFbP�C��W�UMP��z T�Fg�RW[�W�b���Ox��
�6e��픾�u��gdO��`�*]zZ!��:6�� m�b4�vp�.�VԔ�{:F	tRFEoH�o���!
{��ȆT�g@�GQ�}�d�m@�[ZR�p�I�_y�@/��H�dB�O>qN>P����R�
R{��k�������iv���}3 h���O���O!�R,ϐok?4�/���N�I�a�w�w��!����uՠ61N��Ջ�+\�Ň��J|�
��$�p0 І�1S�^�tդ�`h%�9��6g���Ru\��wf�<Qp�:Z���s�|���P	!=��K���@�|֒8����1e��fd�4�/�6�Y0m�v�JSo�l��	~�k�:*�=7=B#	�7��� ��a2IN�1�;hl�Vy�>�9�d��`�[C0�v��{`��6�l���/��ݮ�Բ��"�1jԒt�Y9:#��0R�'�׏�,�U� JqhÈ\��fgG�K�֗�j۟z�
l�p|���!W�`t�V�;Ad�9���� }`U ��K#	��Z�i�0P�dGe-�6��	���z�ŎW��
we�@��a�9i<NH�f�W����	��NH,	����\�X�*\�Q���9��8�����(x�n�ә�]P@U��eɢ6��A�����/��h�"E9�ȶM%�l �4"㾟>dbp<E^�vn��޹���}v�(j;��N2']T'ɩ,�ioX*� �C�:��\z��V+� �7߹�Os��/O7���n�?jb���#˻b�VO���9���}'Mn$�\�M$ w��8@ƥ��Q�ۺs�&���[��4�b��=��Qԁ�$U`���ڃ�)�7G}���⇊�@��tb�0%��]�J�Xk�
Z�z���[v-�,8��t"|�.�Hs��d���W��	dJ>�;f>_��|$������t��]�Yz��GlgVMI��'s�~�p�$��\?��bO��r����!�w(
�� �/��(��ֳzug~N4��1�	Z�� 礳c��O�pR�$,z_t�:2�����~��[VT�F
�B�j�M�E�3HJjYvL��j��
��\ۇ�&f�BF:�q����>�b;QK��$�mMt�Zѷ�Q�S�=K!��w���q�E�5��>��QN��8%Eժ���U~�
�r�%��&��{��\ʲ�1�ܼ�p��u������w��2F��O<�/ �T4q�b%�n$���MT2�h���kA.]�5�Y��؇�zn%H�믠R�M��0V���M�Vb\��-=�X�!�m:\�3.N8K�á+��J�}E&4s������8x�mG�]�_�t���fP�[����5����k"4z@	Ԥ���ȋ��ڎ���a���Y��?����O9͍UQ�3�Nuǩ�v��;���/�_B��l��q螢Y?Ø1��/ͧ���b�m�dç@�^(�ڋ(��7~���>C�"�����TەVArd��ߓ4E��+&��1s)(k�G�'�ݍ�J"��M/�|)�@��®��,���&%�͂E��p�w�[����O�v�,X=������s��p5�H��d;$TL�4�(3�cg^X��5��;H2&_��ܜ�0����>hEG�Xe��d�g�a�8�GM��;5oQ���9l�����2VC�b�k������d^B��a��&,��]15�Ը�����_�ܶ.}��K�7�������$�C� e�E\�^�䨛���y�Dx�8�A�q^AO�}�7���n�%<?�KR?�48G{U�Ov�.�-3�`���������[/*H���A�
�o%)1� a��zgBѿ�&��Mf�G)~",iW�`z;m'-�U�i�����Ai�hAO0�42�L���N�vU�.��OR�Yzݨd? ���9�e�R�!@"��{T��[4\�\�8o}(B\��d"��ok�(��n5,"�fј"�E�����{˘5��I`��j��y:����c��w��#�glR}�bۋ;e��-��P3byTmi���}����t�$p�U��K�mr������Q���{j#g����e/c���4W��^g�b��pA-'y�f6E�T�/�לּ�tkr��f�$D��	��L�/�!5[��w���q�����~�E��y��ka��.��n0s�����_Q��(����Ǚ�KH�	��*��a�7�l��{���Ī`:J�SF�
ύ2��+�L�A�P���x�D� c-=�#?<�H{o"�`�:�t�6�:�QGc%�8�����Q:�������S6AP��y�A�{�XF)�֟L���0m�}WŃ47�����n�x��=�ىӴz�ؗ��,��	Z�UAY��'�y6�BI0a����f���Y�������Ѽ4��vmU*����C�Ap�ɲ�]���y"�
T��F7z�5M}���}� +�)ϥ	������P��_p�G��g����shؚϜH�f�U�T9p���3'�h���C���9,�D@n�e%U�;�7E�ȯD������:K-�%�te����+n�/���O������*�{`�ⱌ���yj񏂗�&���2��[��WR����F�y�Fū����i�qP�6��oUŀ���S�$�-��u�ђ�Щ��4��Y`� �֌���>�=Yo7�r}w�e-4;�m��j�${�[Ѣ���G��7�}����Bv��
����W�$y�4Z���약�R�n�^��t'�/�Ĳz��A_��WB��Բ,��{U��q`�9�}BΛ�8viꤢsn4]8�v.<�i`��>m��x�,�O�J���Z���;˂��4A�U�W��^��igz��֬�@�E����Y�^V-�?E���<RT�)���z��ק{���gAȟW��P�pbDCA9F�J��*��j2��{2��HU3�M�w���|�@�����ffU�9;as#��Q���,ޡ˒�tj�9==�9D��c��p�!��p1�C{���;�$�\�/����BOv��o����nϺ�EKqF\��1�ѻ�}�يMj��z����9|��9���R���Qɕռ%�VqȻ��!��M4�c�V�ￜ��82�:�\-�v}^Ġ`��U[�sQ
s��]�r�ܯ�H���˲�~����d輶G����'�c�e<d�*�3���&`�'�.��q��.bULZ��.�}�D�?Z�a*�ߕ:$����f�U�	jx�w����ܳyy�*�{�;i��䲝�>�����݅b^'��Ȇ4u���TS��3\oa��ž9�'�Z�fd���p�E�Z�mT�2br�e�T)�l���n�{���/6�#o�<l.�>x��@CBn���3��n��
U0p�=~�D�7�_��A�Ϻ�E���jﯧ�Ҳ�ɀ-�⧁��C�[��kS��9Dt��q�Di.�ן�:[���Fь���U!����	����;����<���
'�z1%3[�̉�}ɉ�� �SĹ��6>Ý����b����
 D<=���>�$<���$!S����K짹��Y(˔XZ-��H!Vs�9�Ր�D�ZP� ����Ί%��߼CU���m�~L��(�H�7 
���A6���A��K,Z}�q���[�,�ˌY�ن*A�K�u8�S8�'�U<�L��Z��%2�(M�*�;|��x�T0t��L�����k�quK�I�h��z/��EE����|}� ��'��[�հ	��v�����f�/p�o� �b8��6p�+V\9����A��T�T�i�8�Q4���O��V�h�߷���Oe�j��V��YW�;t�-�
��b ��H�%�0py�c-�dV����<K4=�Ҩ�'Rh8a��j[���r��,���PK�pK���!-���,�Z$O�ub�K���X���k��
��ף�z���� �A��DL�&�G �j#ꎱ��\\ANC큑���kf�(��3����
f]QI