XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� ŝ��y��߷����Ě\���ء5F=L��<�Kk�!	"{V�uo4+���3�P���������CV�*3q�s]D�Í�p9�������A�.J���*���J�zWo�q#��v���k�0��g̈́gODtq�.�٤�|r�[��|zp��!���w�v�mn�bo �x^��-A�Lya Z�u�&WI��o��l\s)id��Sb��O����w���m(��4X��Q�}��R��2 �5���J��u&&q*�����E����굛t8�4��tjU01���R�r����2��|�4_Il�� GpJZO�~�e
FW��a��Q��6(	�ֶ�~����bVfq��B,8d'��L��.��g�7��5թ$��_LƊ\Ә��s���SMJ�g�U��>˔��u�Z�e���d~w�jC��`J>;�P�`{�X|�/�9���D��t:��-����l��6��L#��Z$eq�B�N�ߌ��'"����H�$�v�uTYD(I�=^��ThAfg4�XV�������:��x��1�� ���@���
!rx����}�'���_��'; �X�!_3I�s.�:��@%ǯ_?�#��5	����(g��?��銓 <�w�d=l�+�KcP[���+��[x-m�����(��,OZV�=p��z����v��Nd+3	���ڐ;�����[����o�I{�� ����k-o�*͘1P�\������a/CIO.���<|CF��w����:vG�XlxVHYEB    2442     ab0�%�n�b�'��a����Q���W�$E�p�?c�B}9�Q���tA�*�9��X�V�3�4��	ɜPk��R�DF�.C�8�f�(C���mfq���{6_�/8?�૘��J�2q]^DK��oc�l�K��(�e���p�/���ȼ�������K�#�WJ��C�
� BJJ����/h�s�8w�W&�����~ ����1r�)�C��&�����_Ўu4�\�ɶ�,�:sVCr"�Nv�����x��ٖ#�L;$�d�_	��7Et�:
#�Q/�����iɫ�k��68��w5�G�3 d�bRg�H��,wKJ�����?�;���W�$3Ѝ�~�[�?R/T�mP�P6#�|��g�y#']B��x`�6����D�������b�(qCz(��d������W�P6-�erC�D�z#w[���7[���`�m�U�ih*�Ъ#!l{�v���'�� 7�b0ڰ8�VW��`D�Ⳙ��/��5�!�?�K�.vJ���۱�h�qvEt8J��ԌY2�ElR���T�
.�F���J�ȼ�#4� ����:@��ʫ�ͮ������IC�~�;�_�I��@4�,�M^]t�j�Y�s���3��t�6]��_ǒ�;����@�R��Jr� HOb�8�
X(pF��66�I�ކF�P�G.�J4�XHh��S �|���g��ݝ����!���m������_'��?�6�^,����+��E��ۺDf(�X�e�J��_ԌTnԚy5@�J)�G���©��R4!��P�>Li��b W�g��Q�	�X�E�2�a�p7,㧃�z���ד~��B� ��tb
T&ٓg�>G���87���$з��!��E�1/��1��k0�E��q�ۆQF2�q˳8���>�,����J� .M����9�o�< �o�Z�9��e(�A�?�+X9�b<۟��$k��w ���q����<�oLX��i��6�DLX��d��W�7���T<!H�����f���b;vf�U�,�F=��vL5��	a��9���qv��� �B�����X�+7����������6;�'V�9�Q�y���Z�
��b�r$���:�u���q�ʮw� 熉}0�&�̽���2Τ��gU��t��k~P�IX�/pqU�ů��cFA0���u�/+�4� �]���E+l���8��@�X�����7���c<̧�mC�T.[�|B��-��� �gp���vDFc_�m[�"쇺�O�xo�F)��
'y��&��E9��P��=wY����fK� ��j�c���,����TP?Sx�2�?�sٿ�'N��`�cΦi�����?yA@X[��S<iI��Ь3�0�[��ʷ�@4�j"3i���I�>�)��~��[��mї��D��d��͍'r���8����F�a]p�h�P�-�2�G�D��ń��w�S�#���z�Z�]�䦩�7�����葵If�C�o�"����"�f�5
�#��R�v���ݥ�����
u�����&�M��p��hj���	L+�ɞ��ɝIl�@}҅Jܡ�-����z9�Ќ����{.&��	7s6qQUl:���i�:l;h$�.�![�)�YK� څq�a"*t�oe4%�v�?�I������|�s�5x�;ENH��S�.��l���9��[�v����:l+ھ,������$���m5W��Z �Ҝ��S����%�h�쩛��̍?���Є�3�R�L�dؖ�*�B{��H����2(M���������Gv���7I�}�K�T��D�>�U����CY6�׸1���=�_j?`�t�ɴ��)�/��<��G�	,��,��5�h�ڔ���cb�"M��:
�=��G��S��5�s�El�j��M�5C!t�
�:6�� ah�PYЖ�$�G������3��l�����7�x�h���ֹ��j��x��v�zD���ݘ-	O������1�3��C�����v�I4�	���VXe_�~�L�@Fy�Ǚ4��K�a$��9����MQ�I���������-����b�E�
���Rgw�����EgN�
�!��h��s聉&*����+,�Z^��-�j��,�ˆVǀ�"ڿ4
�����i7bg}T�MS��A�g�r1��t��K2O3��h�x
��}�n��/�����8��U+/ػ��#[��u��s��ֳ��ٓ��T�L����lwm��"�����gV�?Z��%��CŹ��٫���-."6�S^H��\�x�4��"�
.�;BUHlY�j�ް��	$���<��).��L�E����x����L�L���b���`�����+Գ��߫��Z���4maf��/'��uka���s�0�cS�p��4�#�f >��Sc�&$��پ%煃�?+eo��v����f4OW6�t�l�y#��e������^�$�7�w
Q�uE�8�Nr�=�Sx��t���"�"����_�)��|
iA��ȯ�wI�+�f%���񅍑�g��>�߹.��F֗��(n�$*D$ox�sOa�P%H1"r��p����.�Y�>d)RC�A���栙y]%�*��XS�`���͜�n�0��|�P'd:��=�}.~��Y����D