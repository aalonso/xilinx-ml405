XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e'��Y�m���yp�9g�GM�詝����Sɮ�Y�YZ��Έ[򨈎+ߖC��ԕ.���랠H7��� YR�C�#�M�K*��o����r�}��X�ʪ&���[�;�!�y$Al�pʽ�63��.�wr��e�&��&�S���{�	@	��ov�f:����	~�A���0Mb(E�񲣠�VN��C��!-64*��l���W�T��8"h�R�ɭ7���YN#w�@PZ��\�F��L�`��i�M��H����[����B���R� oڭ�|���r��}4��r����]�2�̅܆[�%m�xᇽ��9�o��x��TB�v]dk{Ê�Cw�P��,��y5�S�, z��A�;�n9]B(���:��S��Ӯ|?ɀ��Ń/��j��P�bl@�����h���s���X�092#��&o>��up�1�zLw��u�Jˠb�?�L����ف{�~+m�򤻟ZO�+�x��k_5_����O�pau'D�/L�
�r�n�ȴy�5��p=��b��i@�eBk&�-�\��|���f��s��b	^��E�@���Dv��
6\H|�֦��$l�����ⵦ��N�ʓM8c[��~���S��w}&)tܚ�j�dT�d!^��Ʌ��%ȅ�.Z��u����'O`uc��X�Po�4Yɷ�Z?/í-AU~@!T��ETζ����q:Qt&�A�<�e*�:E/5��N�6�\����y�2�Dp���mg
���k|*t�P�E���^���c�iXlxVHYEB    38a4     d00�{O��W��+A���aр+��H��Ѐ3y���{��,*�ʪ�=��"r�����8C�-����$��a�&=\ ��$D�Uz,��K���
i���g"|�� <�!�Um|����F��Ƒ�Mo�`'��A;�5��8���$c��YCY��6Ǥ�{]I�MJq��x=����ɂ!�Z�M\��@�[� �������P��}��S৊rh�69�p���S�WJ�����Y5���ƶ*��.����c�A�ߌZ��`�q��Q�
�;&[�_j<�{�W*<
|(۳��<<��\.���o�i�iN$%���)�jR�^���_C-HI)�) tg�(̚�*+M�@y�)��f�����b�,=�ZE"s��"Os��1W �Ջ !aDO�pv��*�1Ĵ�Vٜ���倶�M'��1�r������)�G�̍�M�ܤ=���� ���b���ZV7y���LT-��6�\_ҖMЃܕ6�ɽ�8^�z�
G�*����+��u�����ک&��I�'�g+	�Q-�6�����z�U�E�ί6�G�q�|���"̕2
@N�J����D�\|�up�W�=�"ޝ/f57������`��#^)t^�E�v�dw��D)��D`a� �p�1��r#1�I4km�e��q���U���"���N�ڪ���Ge�w��}�Fn.��9�'_��};8��`,8I5���S�ԟ'��h��7�O7�M��D��=B�CIG^aU4�͜�m�h������e!C����Ь-���$�N��K�t�Jj���*��v��%l�?�*c����Sޒ�ڙ�D�L���@
�ЇtX�;�������/���~Gz�,I�	���	��" =����K�e�  ����<�ij(���7��sX=�����i��T�6�2���4�2r���~�w<I�kj�K��^H��#Bז�0�#)[Gl��h�#'Tϔ��.O߾���<s�B%G�S{��^�xF�T�F�Y�9��\�U��N�|����/%ś���ө�(S_���WH�5��?���L[S�/�-����X���H�2�69@�c��o[��ܜ�K�ォ��.[vYH ��j��i-�d�L´l�-��� T�yoNH
%��su�y�y��y]�o�x2ċ�NNzmĬ���n^��mu��18����{
=�����;n�e��'gq�	��4}��e���O������w�\-lZQό(��R&��M�RԄJ
�����������CU,�(�����U�tL�Ao��o;���y	;]2�L��~XƜ|�.n'.`�hy���v���2�΃�:(H�3�&RG/�$-	�Jĩ�����U���Uu�0B���$�x�.���E�C����L���k���<I](C�cx�����m�����!i�o)}vZd��҇�sb_�h{�`Gķ�[r����
F��Ӈ�L�pN��uϧJj�hg@�fXp���?�P+xq�WH j�e)���/�/vjH�_y�[Ov]y�~�Cmx�ׯ���@
��2EV����Q��ڰY�O��(�=����qW�=K�뀔yx���u>h�]=�LSh��颧����pv�EU��7#�gf�g�޳�G�k����?7��^3।�DX�	�	��q��������<�A� ��2��M9�B�"���@�I�r����'�_I�Y p��D���F'2=gB��d����ر��@�~��%8�3�i�7|9�ç�X�2���CR��$u�|7��ɳ�KJ�(�wy��.��锳~dN�u!FH'b�ȼV-�����S�C�������<l����TDq��7�rI��ܿ������� ��F �$ �z�e��}a�+�xc��N�YB�nC�w���qr���6Dg�{l^,�UL�o?:ut�`܅HGmTq��d�L�I��t�=�g�?ғ&H��!_
%�?�)�`�Q�07�m��JN�Ռ#fg���!e�5�#��>J|<[{�f��u!����g�IlA]�cMP;z����H����Ft��%)�+Yn�4��<���<���|�6*X�/x��6~3@����Oة��V�����*���>���C���	]��J��v~VvV$#�#r�T���NЄ�����`Qe�̩���K&jO�� |ʪd���ԧ��Hw�����
�[�i��2P
�d�۔�h<g�<�d�X�o���V���F����jJ�����S��&�<���)�A_���u;�{D�����V�+� {ڗV��05�IVek�?/�V�\d-|����f����}�\_%K�~�c���#���Nh^�$#�*�n-��AP� Z'g��n���쐮��Um��A��쵒��#��YT�S��9d�*�suJ���29��3��+ش�eyc5P�<�nN�Ơ�ZEB9����6C�Ӗe���89}b��Kyo�p�!�n~L�L9���_�	>�g�9u���c��I�tq�0�zF����=�����N	A%�~�rBJ� #��	Ϙ�ឭ��h�#��9�FNb��B�X�����N�&����cr}���j�M�����<�q��7u����2�*c�Xq��J�ooC'K��h�N	S��M��f��*7a��WvP(N!�5��p;�:pD���'�3���$��*の�
�<�7(g��撪A9R�r5�9L%���ow��wSpއh�=>��n�[�+څ&͡&DBs�t��^���Bq�5UT9Ck����R�+��*Y�N^�b}AM����;�C�ާ2��@ei��u�N{�����S�|«:���/ ��5%�9&�QaMB���/�an��{�sX�G��q�\o4�PͰF2�V�A##-�R�H�<��P-p 13�C���L�H��.QK���M}���B���o�(ߓ����@9���g5���ֽ_�'\TՅu?�^�&w8��{�U�"����Vɫ�
m���M���d�A��B�u�H湿p���7�a�uou�ś��&y�|"fQ�;��.�
�����زǢ��[�1ԝ�������M���"�´�n8��];5u�C�-��wݶ�Og|B䮚xY_ua�~�LM�B�Z)�_ C���k)�pPq����]Q1��;�D�bޤ����^�K0���
]�W�.<r�O;FE��3��%�:/��'M"yJ� 6�U�nΰ��f�����$���[(��6n۽J�T��H�/�Z�H%:���KW2Y.b