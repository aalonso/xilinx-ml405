XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������b@P���}��^��j(��`p�$�yt�>�%g�@��\T{P����rԊ|t����H�S�	�Ր��e<}z��k��<Yc����[5��^M��մ�B����ǿY��v�6 ʒ�G:�y�)�
��k�<�6A�4��DY���U�
a�֮:�8j����3��#�^V�6�������YT�H�lN�mW)���!�����ӮU�:Xkc��XE��AWP�ݾ��`���1nJq���~�g�U�,Y�*{� �S&��ޅM�P�U���ԱR��Q<YQ���a%I��� �Aa����8��t�tf�����^45�D�p:�ɁW���,�_��\b��m�R�4��d����2ӟ��c�ҧ���D�߼	}���>���gS�$����S/d�;��D)�K8� ���D��$���� U��x��+"FEc��A��˯������E&�����'�I�:�������5����.�����	e#:ĩi_fL-� ۯ��c�w�A�·~r�T��Z9#69����?���3���6��61n���AH��k)��G�ʯ'�3˪�֯`�L��b_O:��ڪwgw���x�p���}M��k���4�{���<b��X�� /
t�������<B�&��v�
	�Ԛ��"�'�&b�_�:-�r�pXb
-�c2J�;�qK<�e��&�+�?Ը���KV�}P�ԇ��-Z�t�V��!�l)���T�&uy�'��U�ҏ<�(�[XlxVHYEB    5571    1410T����]�C��s(���̣��U� y	�l�oGrb�Gۚ���O�ML�h�QVH�d륵�������8
 ��?�>�*rK3�6t�x`�xGeu��sV�vTi؊��u��p\8\iR�)G�M7�T64��17|�K�ˎ���%��s�x'�?���߭���͔�)�g�j����EY'��X� ҋ�fo��٢�Q,�3s`����G� `�^����u~���wZQM��ns�yh����`��C�.wO�_Җ�t�6���K}�mL�W�����CF���4 O�*P���Gonݘ�m�������|��mИԎR�܁�m�sFK\��l��c(�#�s��1iI|�<���pY9�+���n|U.��0�w�ӳ�����b���4.8��=����˲)�w��)��R��:la�F�Y6�WR��<߃�f�6���Q�����:D�l Z��0۪߭O��e��"O=�d�f��x\-Hfa����pH�B���jf[�X�~��Z��.w����/�jv13����yau	Er�������9��I�6���i�+����K6��9������>�]1���%F��W�H8˷ �}P�_�*�g73�%]ǒ��("�3�֞���"������Ri^�W#P
�#�H�ۙ�c�����[�P����}����u+Q�z>����v7<Q�˭K��j�fԘ���x��,�h��&m�p�$�L!~I�i���22�b�31MX��QJMU�?��#*�'�� �h�xs�?V$���&k�}�5!-:F!��X��^���R{R�
Vg2x�GѠ��#Z�p҆㈙HR�-���V��g�Y��;���d�O��N�S5��X ��IlF5I��Lz�x̢=������EfF����$vo$���V/?Q�[�P�9v�\	�<F�qQgrZ �p�z�Vro-�?��B`�dbE`
2寝@��w�~�Bl�6AG�>净yNACt�sd�V�g�;�b*]�B;ZajC���A8�B{$9c"0��An�� ؾFa<:(nL�����i���q/a��g^I�i�řX��1�T�-ǀ��ej�M'Z��x��'K�ΪSnX��@<V|uW‹
NU��X���\���{����̀�9@�t����BM�EǦ6�x�zr(�\�P;.����Z��d��r�Ϥ=����<R���V����i�{��2�z�����KӺ�6���{݀G��z �"m�	����jc�U��?��̾:�5�NA�V�4����l�N?HnEpl�rT�O)�:�?�eV��AS�-�[<Rj"Z�/��L��7�uZ�M[�t��g�Y�T�6!ȍ���W�Y�M%��,|lP���e5H�v�4��:y�P���l�O�ޣ�i���*w:${	Xx�;0���l�؎*�5���~ľo"'d�����Â�̼)�j��:��3��GPf��'�@X.���3^O0.���(��яY�~[�k��%�g�:��C��2��[g&񶻦)����j�4Q@�K�'��-�$R/j�@=����/�k�
�7@����Z-Ox糮�_�[��S�-�� 6�ky~FhA���էL���m�P�4����SGiե�-w�� �К��֡P@ې�U\~���_�5��jN�Յ��C�Q	ݖ�9Q���l�2jyǕ����_�}������Sԛs�������ٱ�l���1A�C�X��O�)#�C\��W���:�M��+SjEL�����s��ȟ#.�w�M��k�4E�'���
<2��-�vn�N�!W-7~��׿�x>��@Spj�ׅ�1
b�����5��w����=�����(=��a���Ld��9��LبʾDd�|X|.��+�����c%a�"�~���=o	C�G��-���~TUEʞ��X�=s��aX��ó;�6��� �E~#��zʓ��k�E?E�`TgҎ�+���@"A4����a�i�b;m�	
�,F	�k�bַf��.�E8���GA癿�L^�"
W^�5Xig�+}
\I��,�O�:�P���eHdO�cγ�Jӏ&�'Jo� Q�iYN�s\�Z�� ^�r˼l������@�E�k��>�=^�mN��UpG�G���y����G��gN���((M��H���LҾҾl���=l��I~�,�1�T�[�h�tU%^�= W)�vB��f�+*K��c	ɂђ�)k�_~�Z^Jv�j?y�l��YW�U��9���Թ~"npf��1��2R@{H�/KTOx�Z$'5��3��<wN����km�%m�a\�yn�l~��0�D�� ��n�-��I�����(�����wnJ�!_קա��/u�E,�����w|y mx�/�T+�Ym�yF���-�W0-]������M5��	r3�;K�t����5����k�`��Kcbr[PW��w��K/����Q�������8;��ɻmF~�tN����Fq(�/Z�ٻ���j���:���N;�d�K�G���n`��j ���@z��qO`4#
(n0̮d`'��y ��I9��36u���o�޻������{SR�0��Ą\oX���Z���#��H��DNeh~����*�9�f��k���{�(���ǋZ�46����cg��b�O)@��v�����X�r򯋝rq�o\�g��n�Z|�ze���d��(Hx��8NY\y�?���H=s�k+���HJ݁�J�hR�����-�h7W�'|_(�Z4g�f��"rb\{�u:gι>m����Cb�]�v�t�M�X (��d�� +�3���E�{�	#�
�0�G���${(˙�^;5�֢`���������w�����Y!��>wL���'IIv�#�R���=@�J��;�Mo�|E8T�,�ɯ�ɲ���^������JV�򌞌����N"���8舮)U��{�i�9Oh?i�J�K�q��8-��c01���{v����Iz������A��fw�@!��:!p@
�j)__�A�F|b�-�S��SU���+�J 4U�\.�EGa=h��c-�ox�a��xWR�Di</�A��&�<֫ܘ+�<�h���5WM�1�\�����>�T�ș.��%I1Բy�7�j<U�E^��r/�M���j< '�<<����L���UWZb& ��s�����k�f��P�4c�:��t$~��Z���9K�����u�r;O��P����=�{c����s��.��;��o�ˣ9�E���p�ynRP�c���
/����r[��G'��3e������A�����#�6z��q�ºy�&��ݠ�=�<rO?�ThѠP�l��TſY��N���te���k1�����hhc�bOA=�4Y�|Pc�l�?�l����{�D�]U�5���\�R�c������m�����Y�7�D~{�'�s���S ̿�xSVM�K�}��b����n#w&{Ux6�a�f�!��o�����tc	g�x f��*������f�S͊��8��6���u4�ajwP)��ji�It˷�����#*��A�]�@�2���ԙ�"XsS0�9��'���q����62�(M����f���Fw�x��hM�� bMs+*�TK�5�N�,�W�;�U�:~W����<��վ�kV$l�=w��� �ͷ�)*��NOD��}8���=����<}q�� w�,��e���@F�b��Kv���"�x�`x��h���w'��f�y�"��(��D�>F���i+��Zжo�_k[i�J�J��$ZP	��,݆ N{f�e��>B�E��<��8H�kC�N��6!Z#��J�Rd�&+�@�\j�mG���������"��si�~,�J(�p�i�#w�� 9Q�7\Eڂ]�{��WH���{�����p�� xe,��,��ݴI�yW�+�X��r�#2�sg��s�b4?�/�N��-�a�7�Z�<+��
���"7@�*0[��*Ax�dL�����j�]��R�"c���7hT��c%nk#W2a����l��)�����gtR|&���x�'�x���d�_Z�{�K�;uzbR8��{�8��-5�+���c��lH�1��c0� �'�G���q�_e"뜇ՃǢ팑M�i��X�O�e?�O��]Q V��Q��ڊd�;5Zk�����r/|3,[m2R�L,�]��ΞS
~G�K� �� ����>���јHq�%�!E"��x����Z=��$8 X\���?7���/�s�s{IG��:J�5V�[��Zv�d���?�N��%o�8Kjj܋�W�F$����E�v�7�r��t���)Jx�}���S� H�ABD-���TQ�=K�V4E~opi��,P�d�}���T��i~�fsq�^_i��6��-�P�_���������m�d��}c�e���8�Kz`���F$:��X�si�n��)�1:l	� ���.��]�GvjWO��K�����e���z���uEcz����~��A���A�ԛ0Q��\4C0k�.���qi�������ǃZ�c�}Gԉ`
�DJ����}J�����!e(ópa��+�Aљ�47��(}���=�"q��H�?b���}_a8���	w�ᘖ���p���𞻋%��|��-h��"w��A�#~��]#��^aQ��ܦH�����4��Zt�h7&R4�?���"Ϲ�3�������>��袺-,ω��.���I�"v�[Ve]=2����ݘ��Ȕ�L|&':� ���.��-мQv�8����)���B�e ߤ�D���T��Xf=J2���dB2!����ަ��x�(�w���d�K5#Q����y�(�����7?|�dT��.��1Q��*utjF��.Oq���s}]���O��������Nhw�&o��b��LC'2�n��L�`�����|	y���O��+���g�v�F'�zb�U.�}W��^���1E��l�i���Y7r��$��r�0�ЦYf�v�pu�P.�ݰv��D���f*�Ql+1�%j[Z㑔�(Z�w�WK1ռo7v��0����