XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��J@���[07~�m�}���}E���9G���Bdd06�"����y��.����y��-ѐͪ ��\L�*EA��*��#쒝��H�s6N�6��;���x�T]G�נhN�����H>��{�p)w�0-���<%���bұ,�&�4�)�����&��qT�CB�-�K@w[q�r�Ə��3?�+#%��@� e�Aj���Yt�w��+n�^����l�wjO&G�'��M}��z���饹��_m�lh��ӛ��#�-��r�O�t2�K��mz��!7�&*z�Wj�X�:=��������)�Ă�S��_���m�]��k���s�9�h��J_���x/��v�Fz���gbH��7�����̐�x~]na$@�`�׍=�W�̗�sK����>���@]b��ފ��k��	{��4@B"�` {�p��{�3��(~-@�����sn/����v�E /οʉO���l��:�̐��I�N�_�E�%-@�%�#���$'x�ԑ.�jc��*wA��S,2m������n�lQD�J�8���y1�sD�"]�0��H9���7�<uޏ_�[�����3��j�ȵ׍۩�38(�l � ���*���O^������2?���Թ6K��z��ED��R��Z�a��ρi:2M��)��n�%�j�ȇ�m�2����H�x**ZO�zT�כ��f74��>df�����ִ��{��W�	��z�%C9� 0 ��~���]�;��k$�����70�w� f"XlxVHYEB    fa00    2c50�
�Khtk��/�2a����� ��!���6������`m����Y%W�4��N7����abJe��C7�S�43�$o�ec����4l�o�,rv�D�2��Bp�o��3A��d����I���B3��<*�:�HJ�e՗V�
Oң��@4��X��{�/p��M�s�E]>X^b��,Ƌ(c0�@�=�O\.[ǆW�qJ��q�}a���%T��d�z,�n����K+26�r�V��z��,cb#5os������0�Q���LE��Ä�5��^�8ۀ�g5ڮ^��o�h$�`�׹����]
3Qs1�>��CV��	H	32Ԑ�'�b�����f͗����M���s?�د.��{أ+�,�6�)O.�4�؀�����GU�
�.��-�1��Osi�Ne�'�L�b�8���`��{T��N׎����.��/Q�H��F1A���̘m?s֒�sG�αW���F��#]v��m*�1��k����X��n�D�$Hײ�RMV۴7�t��{�|Y���'�3��T��&E�e�-㓵��{�l)��E����i�t�3���w�*Z&z�0�����y
�K! 2��X�4�"�w�[�4XJ��>!�K���2P�A����s�ἦ0��[�湶O�b�R�^��~��_PK,~���;Zq���(=Be��1������#���+�&�[�Gp�qu飲��6Afmc[BB:Y�A"V팣��͌���'�%�r�e�fho�Y�W6d�kF욛y���䘳��3�dr�<������J���L긜4]���!W~�q�p�;vò��cr/��"yKT}F� �q�i�MM{�<���cq0-�[+`���J�KD���chb#���"�ރSuV(�o$�����6l��#M A�Go�Omj���\�]���Ox4�XT�H7�h�0G,��v��{3���:����7����|2*�5a8t�:E����a����)�b�뉇~��7�%ǛR��7Q1'�W&(J)O6fTc��1P�	�j��gp9-��j�P�2�9�=j�V�(����m���~o/�;�Ԕ�%��V^x�[�F�� ��Z�8�Z@�<�(� �(RՓ�㐧Wy N^�VN�X�p*/s��J(�SόvU�ƀ����[�b�M����H-m���=��	�3�i�౶n������ ځ���μ�H0�a�G��`'�&�T|-��p�P�uo}E�r{��֊{J���/�_��	��y�[���^�z�?�?�ضO*��޿�p��T�3\1z��=$d[�{y����1ތKP�e:>vH��[���Q&Q>����m	�8���f:Tʘ�3ikgS
~�]��(�X���tc��)v�Ks��-��lJ��ú�"��q^dN	��J��Ss��]-��T�UPe�ݮj�r1� Q�E��	L4ܜB�����Y�1� ��}b*�m��˪C�VsEk�!k�b�d�&F���õ��ѐ緲�\3blr���u�A�i�DS��ſ��}$�N�a���ٯ�U
q��E�D����Q�J���uN�E_E�����9"#�p1I���v���1	��ʭt���٨g�����hR����
�⥽��7pܾ9�=�d�*܆���=u9˨�P����@c�3~*vc_n�E?.���|��u@��nwr<����ᇅRn�^i9��ߛ��U�m=W�%�(�~?v�GnN6_Իj��R&���Uh���C6���V���M��.��cgi�o/ם��V����<o.͎C?N}�!�Z*(���Wn@l]�R������LIp)���'~F���gG�ʖ��7Z0�����Y~�㺼�f��lî]@�-`��Rڈ�[zw=�Ũ��0ѷ5_`N>K�,zԗ����+�ei�	�a"ռ<�Qtdq���f]��&��p[n�E��]�j?��<����^lax��&9y��~��x�6�Vn�hd��?��6��N���G�;��v���]?���Z�sZ|OS�-��T�d>X��!.�CM�H\o�x��H�����R�B��J!U_%;�~j�r�7D�ʝ�j�N6ss�����b�kʶޓ�L�N~~X~���W�iĎ�<��~�@�V7��Ȏ������ܤ���o�3�D�#C�ʔ��'̐@����irI����4��{�)�.q���S��|�6QI?���:z����
f�2l����p)��w���~	�sY�r�:�1��Ѹ����f�,1�b㈾ٲ��h�I�g�rⶐPs�]}��rj����� �?]�/úQ/�@��Qsk&wNH��7eS[�і��j�	х ���a*}��A1�i�!8P�� 1����~��EH�#J�Z��iK�#]������]��8������
���~8T �U��,�b%�������M��	���޽Gƴ-< Rތ1B���0�M�PQ�u���O�6��Yi:/�����'�o��hއ�i��2�?qI��֤�m�,��r�|�D��RF{�'չ���V��rL�3�R�p�3�� ��v��!�:��$q�̈́�G;�^��!�M����d1%p�
��|/{��u"e�(��e(݀�X�jڨq��f��Z�P�M��u^�f;�n�Ć�B�Y��6قׯg�v��.0\�����Ӓ��&fe7LP�"mf7�¾}�~�!�9Wc�[=���\�+{|�q�}A�G\�U�gf/���NTh�QL}7����9�砌�#<�^,b~���ď��dZ�p�e��	��x�]��	A�AaeG�;zL��Q�7�k�d霒�uGp$Iu��'��3��}2��zJ�^���/Ə�:-q}'�ئ���8i�:*]1�6���>s���e���c�={?K��B���J���Q?[I��f+l�N�{~��n�~��{a�E�ð��Fg[��k���%'���v����Mަ���=Q�@8���Z\�~?�$�u^/�/��nKѯv��?�-Y&D3���\�����Q�,G�gJ��f��©���6�H��z1� {Dƍz���DFW�H�k�"4$�K 9V��R�)���׶Ke���}�MJ�e�8�uT�ee!�6!DB�u5����#�@Dڬ��F�L���5�Ѧ�]q�5Ty�Ƴ8R�i���Y�p��:W[����YYܟ�]o�Ũ������~����=��	�R,':�����j���z$0j��vEJ&�1�����N�����c�-X!#�m�����0�\hX��!��C�pI��n�*
b��<"Y��;hܜ����%�@(\;^���v%O��a����	C#؀�Sa�5��S3$]�?�L�ֆ�sr�ڄ�2�C	}�Z�ȏ&�C�!����􇲇;���T޴�#c��z[��}�]l����Җ\�otMn�j�[��� �!V� ��=^}�p<w}�u�<c�Z�����P�K)a�4z��|c�tH���C�^ۉ^/�4Wa�m�<߼Ni���nz�G�Ʊ��/�Ȫ�މ{	�R�Ÿ�N]J4�\�]�{���3��-���{��kQ���N���O*�%u8��DՎ�KrL��{��
�]���%C�aKF�1��/�ļ%�phw�x��l��ؽO|2�����hIb
jM�����Ԙu����N���IMa��9|M�^_*0e]Z��{�vܞ��B�$���G�I8 3d�e:~�A�8,�&��]�*���n���_���̡j��\ɭ3`�J�,��q��7�W�N"v�
��[����kB-Ț?�D�p�o$i!�Fݗmd���7�C&��eA��!�gh��*.V-L	�Փ�!��"s	U���f�'������]̿�I!0�T�A�O�w;�(B�;��S�L�W�S^7�.�)�[88A=K4;���SI��~�oe�?�Ѭ ���n�����Y&���1�H�O���g�p_U�IRC�N ��"����$Fe�����G��(�W��j����r��1Q%d+���8��h��ssf5�eʔv=]�)j	w����S��l3���� �N�>iFô��V0Wӆ4�gV`�9��|Ģ��e�us?�� R�����9�c`�����In��,T�Y��f��>~ڳY;�+�]��
F�y怂7��ܞ>��Uk����5�:y9hh~��B:>q&�;1�A;��=yh��&93�I�9�2P��ą��H�$���0$��n�2����R=(s�(��R��K�V~������ts��6Oq�F���^�������s'���W����{��k� a��|�Pm�i8!�0�5H�z3��y�������,=pe��� ӻ�����]@h�F4N~?7_[�
�=�.��X ��g�\v��K�X}ĕ��W�=�1�笘�c�����̌ˤ	��*�bE������
(!�>l{��V�f���I��7�V���ʃ߿�������T�hI�d�e�$B�엝���H`���){o��O�*v�}2��L�0��'?YO ߯�c�P4X�V�����(?�q��	�L�%B>��jWU�[ŝ�ج�]"�D�:�AJ�F�|�H(e$q+��C�9G�G��_'M�}�%�M?�1��5n~�9�U˭��"��|�<���x���}���DkY��k]��ng�7&2Lʷz�D�:��B,}���/-U���C�_��a%�t*+�Q�lO��wE��F~^<���Z��������(�^�/�J���CIz�$�AL�X	<$S�S�O����+��@�̶�{Ŷ[�'.w�|���ϕ��ތEd,,M��O
�.jA��Q���Af���DhI�e�B�|�e"j\uBf���n��.3��B�6Tbl9�>j�k��>�֓o[�H�m/ܓ���3<or��d۳>!��] �ع�jeІa)���ʿG�����"���s�u��h��o=��B������ D��I��_��F��e��x��@8*S7��������}!2):�ɹ	�vx���dOìf7��yWk�;�{�����$0�ʳj�y������o����Zm��XB̺���K�����ѕ��(&���}�z��mՠ>H���&*!�r����(���lՌ��{MGO�^���%�k�Ki��*"�{����(�x��֤�%<�Sd���چ��v�~!������A�_M~2L2ZJ�}F���E�4�+�e�L��  ���=,��s����s(���
�i�|��N�~Q�/D��5_X�H��옫��b�yCP�I&��w�����%I򉚐L����K����lj�0)d�{mH/Eh')�r/�3�l�6[&�2�&�r�u�ij�/i�I�p��w
]�����Y�+)-���L\�񿢚����AmV�&����އ��+��iB���0�R�ja�Q�ʽP�(b,C
�����`�O��fS�l�N�9���ͬ�����J��y����(}{Eo�j*�%v�z���6�m�[�)�s�C���Թ�0��@ O�$u�s��-�E�O�P1'wZ��lN!�k������^?�z�D!e]��#!�7��S�R7v�?�/C�a��Y�,�뱒7�T��Ϝ�(%�oz˦H?P~�?�lDZ��;������&c���SXJ��r7V��*�\ww�W�i�nR��J���x�|޳����*��f����ED���}�&)�$&Ap9�� �c�Z�:�u�O0朔%Krj<ⱨRN=voG�3$4�<�(W���l"%�[� ��e�P��>���} ��3Ϯ	��N�zϙ����\d�)"x؅��?6��:�R-����P��1�g ݸC���(a�o>�;�K?J@00��ӑ�?���<�����eS+m}g��13�&W�o3��u�Uꨴg;ʿp�R~��>2s�
��K�?��q�� �r����������,�^���y�wQE���M�Ķ�+4��߾iJ�	���URS���o!Ȳ!֠ΰ9�w ���Ѱ�y�^���c��w��8[�Op�t7lz��PP!F���~|�q����2ͻ����9�;J]!}�6�Y*��ڻ#�� ��2z<�����7yY"gB@-*��ZH�\�!l�إ��n���� T��G�C<��)،�����^�@?7�i%#�E���陒Ŗ�z�֎��2�cw>��ei�ip�G��ohLV�Y��YI�;mi [��ȻEm�-eGId��"&�n�}�
�cl�۞1f
ڣ�&i��bj`��}���<Ă����^���j'5U��~�s�JY�?��6�e�>0�����y�۽���=`���_��i��� E8/=X�'��n��܆ѣ8cT4��0�5���Л@GxR}����#�N��ԝ�{;R�P?N��d��6E�!634#� �]^�_����`&��s�q�ğE��$"�F�J�ژX�Ю>)_�2B��A$��ƌ@t�� �&C 4�Ȇڛ��	���@�>v`I��y��{�=���؇�|h�5Z�L�5����;�-�qL[,����TC�G� 7�I�V�J�:��1�΄����g��
�����i�B�?jǋ�I#-����>��'���d�R&����M�1ylG�o{�eA�:�^�i��x}�m��4N F�7O9�!�Al�M�o�U�A�<��"���f[I�qmM�
��4�c����F#7�{D����X���ʨ�8T�C��嘮
E?���>R�Auî~_M���wй?�"�EvU4-yT;hO�Ǭ����1�⊴��P�mr�#X�4��̩�aR�(�{��B��p[}z~��L1��F�@3Ѽ�MV�J�Vl��W����,���Gr�k2����0��Xd�����g&�h��2^�n�k)�J�Y%'����a��K����9��2��8�+)P��&I�\7�t�Z6����dbk	�.�Mv�RJ��`'���<�`+��w\B�x�;�#���h��X�XI�i��mb�.�UD�?�B��O�n
r�.T��
1�)\Q�]����竐;H){�u�Y'��,��00z�p �E��V�bՖhh�Ҧ�׶���!�����-�/-�d<�q<���1����z��U��	�(��i�҆ =h��	 g5H{���:rr���� >����ࠆs�� u|��΋<R\�;���)���7>@�2u�&l���&���#���^�3v�C'lw��B��	��B !G3_1����,Pe�C���&pQ°e��e=���[�Ke=�����!sܑ�Y�@������B�j�E6�[���cT�i4�@[��p?�@~\�� �V��xYe+�|4|���q&3�`!B j9�dq��b��d��R"g���V\~�ů;�_�Y�џ�8�'G2Z<Q���C���i�e�9�Ѻ�_π���;9�X��3�E(x��ڔ�nB�CLE�Jِ��q܏В�h��'hj )?/��|�qb�?���O�u*�5}8�?���j!#ӊBV�9:�WW0������ŋb$q6S������p���9�p��I��@�z=���b��iv�3����KG����b�S�9KT�&��'�FJ��k� ��-�{k�>Vk�p��B�-��7h�A���u �j��7@WA�L6���Q�nBm���T!��[D�aއ�]=����A����]4���4���3`*\�>h��6Via��=���ye*jq���vIlaŶ�yԘQkڧ��Z� L����p@� <�1���
P(�|�޴�0^������<"A��6]ٳ�7?��P&�,���w�B�(�]#��3��4L-N��N����w���q[ͱ����	�&2"��o�O�G�.�X.dXL%��-�`��٠��lk;'lMV'5fx����@��[rs0�[������k2�ث�?�ry����mE���&���~�*D�3����ě��^�L����(�s����*�;�2A4Y���xNH����6����(���3�ؕ�Q'y��:�?1��mHbp1[���	!X�+���6�����x��[G���˂�����o\l��	Lp�q�43�k1Uc�L��w2�^��/HX�<��D}7f'G���:��l;�U�����s�k�O�wC��uȧ�VїZD���$<PL��8s^<�8$� �2#����"rWG)Ot��Uq <t׎'�-�?��HIɚ�0)J�h�o�+�3!��
�$��@Ü�hj�+fH�C`�T2�wF���q=�opls��j۝	���f���2h��{<Ն^���5��SQ���u/�ta�/�FM6���%;�k�=�~pw/Pr��*6��J��a��e�׹]Ƙe�wR��uG�{r��A`=Ʈ�]�	�sHnF�%�:)���I<�.������� ���f��u�BT8�x!M&Rq�U��]��$����<��o�:������'�I֗A}C)����;��U�{��9�}u�}���x։��l��k��:�>c�Y��@�C���ϽMb.�AOO���Zh^Qۼ��v�ˉk�����qꯝ�����v�|�iT#������J|�
�n|F��\�OV1�O�F��o�vAK`����mg�,ŏ@?�
Q���M�ψj
&��r��պ�1��!ںG�<���5Ī��4�N9�{q�1*r��]{=�Ll�	r�{��_w��c��h ]��A^���uZ���n� ���
��c|+�!��/#rOFn;L�cˆ�u6���1/���V������N[����H�Q���Q�-Hc��qAc�-�=a�5�ރ���*������s���TҀ���9I�ƚ�'4��be�9k�k�-��.˝���oF~K�#7yu\�I���/�5!�n�fƯ	)�J��BUd�гK�i�6�9��%�ɞ���u�>ѕ�j�˛�ǥ+�+�j��Ď�ҹ����6������Y���4!���Ь��a��%�T逯��P_�:��_�<1V��S��$ѳ���b~�2�`��T�s���N9�C��B>Igu\%�)?���4�,FA���S�q�L-
Xp���O3�S��X�Nh���L����,"I�,����0Ũ���_g%6=�{@����-����3�k&2���'��D77��6U�R�!�	/��	"m��mH
N%�
czL.,G��+�Mau�WZ�$R����L��]��^Ү{�##�a-alCV�j�'��p�'Ca[oP:���[�]���-�`�e�����b�(��1���d�In�E߷���_��V��̻���&�a�أ�;o��'
�!o�3rV	F�GYH��E=�1��&�|xs�gѧt�}��o�cX��̱�=��E��5��HL+p~g����*�<�!9�QT\�@=hH�)[e�{I-v�8��0˾+��K�y���x��f�Ń��3�:�#}|z7$'����,%�!��a�T���A+����B�~.NP�@ڶ("u;�n�B� �`�Y��M�J�uK�Q��uT��C'��|yv�����m��X�����91p�i�3�qq��E&��x����e����R_�[���B7Ã gN��F�m�lE�Ǐ��,�ݎ�~"����7��C
�\�ԿA�!q��|M�7O�Uv^r�Un��Ӊ���=:����9;���+�q'��]���3�'�Z�̄pX�`���Ψ3s�E�< " 3��Ҟ�~C�(m=�/B5����j�|��@ �PI#��{(	k�HY9�f�W�O)�2��F�>�5W�W�R�}�S�VI2T!0�輦f��e|IF��#&	���^>e�}D�.� _��c���-�������� ��E��U�����r.N{���|W��qRfZ;(~wFx�e�F�|����/��f�\�˘ؠ�=����3:��P�i���B�-��%��{�F����iۚ���$�b/-|���)���N):A��-#��2���97��eo-�)�5;%N�4|F_�I�X�jz�R�F�5���Ba���bep�CһY�j��J�_�sؐ@D�x��{��myb��P�{KY4��r>�o[Asu�AUmU�AZlh�¤(Fr��rd~G����0�hy�$KW�5A�4�oD�ޔo�)hK���rA�,N�`#n��Ou���Q�Z��ة���s�w��"��������&鳮	�Ԕ_{���l�r=�AU�5��G�Gԟ'����T<�s�5����p/��'������#�.pu2o4x�~f!Q-��B��&:��^����?��U���zKw��U�Y��q�o9��,���{�����?d�߄�2Z�Fߙe3A#��R�p��h�9�]+���P�L(�3�C��|)��Մ�D��Vͧ��	-���n�i^��OgY�c�4�XU?k�?>gE!i�F�qp��5A[�І��cH��Ck]�6����5�,hdtj�/��bH"~
W������nP��$!���si��`�|�i�=��l��{;Gؕ��DMy2��
�A3�|�<Z9sC&Ʈ/_`�a$��x�2�K0�����/x)�zF�	�k��c���:b�!#@�?$�"�q>���ՋЬ��E��|=�۵������taz	Z�6�o�x���\Im����Q@h�<�+E�R����w���U�i<1O��1ts��'D�.Ť�����Y�l?��솽ɖ')7���@c3��R�\,��Te���E�������sb�f�F�f�zX�g��e����Blf��}g�:�f�+C�fx^��{`� x�$ȏ�9	�Qc: s��ZW�/��[; ��؞����UN�J�lH�h��e���Cx;�uH��r&����F����Ѷ,L��'�E8^������R�\��C�G\�z�T�*1Ge>�D��6�8��)��r��V���%:톈���i�v����*zYLъ'�8P�xS(wǶ7���`��*������S���l�wPO��ҟkR�z�
g���Z�?�c��Y�UĂ:�J�Q��6�a�L�Cs^���l0�d���S:�um֤���
L�G����C�`R9���7h�Vb�V�?��O�;���D},�}8��$"��_��<�ź�0��M��r�הc�cr���DO;*�mͤc)�\�`XlxVHYEB    c397    2030I�r����0]��XZ�}��G[�v.�G6�4z� ��`
���yW�o�w�OE�����G�G�ndn�{b��lק=�6�|B�丨i>u�I0�s'�����ϼ�h��X�����u+c�1%�"��,��q���{_u��G�Db��B�P�z ~d�ֵ��b~���u����kr��ʹbd�v��C�y��)� (Z'j�kE�ɷ;��h���f����6_=u�O�������q`��wPְ��n^z1+�\�c#���3�KE����O��f��C|P!����-8H?\=_r��(�TNA�p�!)8����<E'�����t(f���������׋�jȞ_�X�K;w�sd�˜���(���x�'e-Nج�aMxO/K�!�	Q�rhn	�C�@7��0�� �π���sxz�J������>��I[��3h�ն*]h�d�]����O<{�l�i2���k(ԇ"Y-S��~���-S�W6~N�o��vh���#Cu%��H�� �l��ג�y��ad[;���l��!\v�֠5k�s��a3mYENL�9_@W�{I�,��6��0����4������W���@�}������N�	9e8�sgd\se���މ�7՛�Uu�؟ ^�<�&�C\��0[#�x� � c���e�>Å-9u�ڌT�0/��{�Gf9r��+:�?�9��R^��p�&�82j"���u�5���1I\�I%qפm�o�s�GS?z�ӣ��0�\I$��6L��T	&�8F��mq��X���鬘�I�݄����X
w�P�yf	�~`χ]� qܨC鵇)S�`h�e��=�Ew���%��Ҳ�D������&�X��CU%�h��bt"��w�c%����[謖k��\7�.���Z��,5��CՁ��&<�Ԋ�#��7���3�a\�U��]pK�  �򮗗�|�~�P̮H�æ\$Nn`��%���l7jW��$C���y�ѷ�(CLd���N�N���(�btÝ�0���}XE���1�:�p)����&ݙ���>Q����_���,������3[�@�ω�vb�MmN|�����>�I�4�dB�^�I�J!BO+���&쒒D�6�Pn9�ToN��X䅨	̸��3�^F~ŌhE���E]�����c! �0���܅���o���KP^�$  ��T\���@�I�e?$�X_Y�_�T�Y��Ë��1����d�m�)�k�����D��67+7��F��/mqQJ��ÊB!�o%����ڵx����u|���-`1Ќݵ�x�
��i�;�t(4�m��'�(��!���t����C�i�6�PF���T5XK����%z�ik�Z�n��ej�n���&J��x,h�T@&�"����<H �������kDy�������:��`�1�2`��{̹p�}�Z���4���T����	���3�c�0�^���#��8�fN1~��������d�/��:�J�U0_�X@9N�u��7�-���4D��0���R��>�यT����N)��	C8�i�%Eӫ�{@&X�������f��
��[k���>F\��c���+Ӌ{��a�J�����u�+�e�"��d:�h��~�Ü�t�L]]3z|�B��ʣ벨l�+�wfS�H�S����>�j0L㱎l��u;���q~�������E���T]Y����6���u+җ���q$5U.LZZgQ����m��$��b��lY�@I�.�i�aM��TI +$0�Ee�������l�O�yF�~/c��VDּ"��R;��]�qָ\]Vh�k����b7T�$�۴�忋wQ�C.��ٞ@C�$�uU�t�`g�oF�8;/���&��q�h���̤�ܞ��C/X�!��3��r�&�Xvۣ�V�2�eT���D���F'� A��@��H������aG�{cX"X��Er���o���6��r�4j��?�<���ۜ{�3:p�_���EHoI�|�f��0�S�3Lq|Z�]���C��BV��x�6�4���Uޯ�ֽj��!��E�A8����&w\@��H���|�Je��L���L�!��B|����5(̉�P9��-��P	:���K�V��{�,SҠ,�Vr�W�MuR�U3J.	�qS꓾�����ߘh�I"��B2���F� BP>99�l���K+�j�,6(���qGN,���oK4���V�d����\�>�k�Է�@�j��i�4(?Ʀ|�Ĺ��d|���C&R�8?9΄	�)5��CM�*��
�>�ɂН��X2B��S�k	=�<��]	�>Ma(���,XGz*�;��`Bx#q��:.�%�K�k����'����U��]Ý$ݵ{�]��̦�0u�����5� �p��3�B"�:���i�o��P���]�zb��
?�vy��U�����\͂t����R�1����+r}?��r`�t�L�aP:Ƴ>��q�w�e7	�.�t3��M����q�^Ú����ݕ�@����a�τ�P�gYy{�l��[����=u%���ÚM fkUy-/���ݔ��q�R����͟�Y�Z;����J�4k	ȟX�nX�d����7R=�T�O-��!ڪmP9�ht56�H)��كV���67$h���T2�|"�y/2;�q�\� t���_k`�&��:�Ғ��6�0��nu��)����?�t�j! �7�-{��&��&l�R�[�������c]���/�!����F�/&������@�G*�~Q���2]��z&�ȹ��j���k�t��6��bhe��D#Ր0�%(�싔TK���ꋮ��U��(1OcY*���/�@+�˻B�9�or'k����e)	8^MuƘ�O�O5��\�a�ݪz �Y{ hN"Z�
����D%g��P�C[O��[H]�E�b�a�ԫ/g�q��=%N���.���WrAOV�D�'��H�o�]�Z%�� C/��>Wd5�hq���j����"%�F��P��{}�G�es�I��ֲ��>����m:w,�q��W]��C:]��sT�#S�
n(�ڳ(��;���fJx}^e������>鳥&�d^Q����)�rĉ�wI�\N�W�U=����ɵ�m�JhU�8:Gb�v�E��xS���^Lb#E���"Br�Xm���֣�6	�%�bhAy��^���%ݛ�cU�>��.=��|�����\S�б4���4g�D-](��:�]��6�v�C`�r�W��}5��:An�6d��K}
�1��U���r�����וz2�"0}#R���q<Ea�kb�m����u]z�Dq�*,���nߗ��>�[ڠ�N� ��K�ѽ�8k<ߑ�p�bO`�8�q=�|�D��5�����4x&�p�۳�o}|�+;1���8?��G b�F��)�����߷�yQl�(�o�r�n-{і�- �o��3-�=O��+�D��E.�s�%J�dՒ�	�ԏ�jP�0����� �[�em��y�cfy4@u�g�{n��#] =��ۗ��0�J�̦���-L-�l���]���z!
'l5�z���m?~�R��#��Vr�a��]T/��Вoi��I��P�O]3�z�*g0��Lx�H�^D��Ry˟�����ңZ%^UUxs��8�%���
�N��6�>�]��9h��n���=m�{��A�h���8ϧ�Vu��L�W�z��+��RZ��=��o�VKmb�(���R&4�z�kҬ�G'gI;?D1���:.�N/�8Y����^fa%��G-ݓ�{�8��jY(c/�P�[�Tl�p�a+KW�X�_t��j����Qc�?���=O��� /g�zO���r�.��o���t�ky<���T&���6�t4>!e���28MX�X���R�˅�5�c&{x��?/nT9hwf��
��a���������D��J�f�km)Ya+��l��>
X�TONL�-�~���$4DQ�g�~��_N�+%J�BB��lR1%�;_�F0�� �t>n`�����Sܪt�zMr�aɹ�b����p�C`\�	��twIw~�dq{�_��*$+Ԕ�;G�Hr��7�n�	þ)Qb1f* I�É��8�.��Iϲ�}����y�?e�T��oIlr�1����g�g��s�c��܊h�:DV".@�g�����Ji�~Xf��Jr����Sv��%m��
��,,���%�W�e`gG���P��u�Y�ٰUg���1��1%�J���՞޴�ב��g@IY�=ha�P��^"��9!�d ^K	�3@��8\_~!4���v���"�����*;�R��s2,�^�0G(�a�x�gյ.�{(�z h|��t<g+(���,�Ď�k�?��� �	�hN���6��:'��,�4p���Qto(�P��K�9^��Ċ���uU��w~C&Y3հ�}�V2E�-6��+_^G�ȱH��L��jG�?��e��$b�Nf\���r��.���6�"��a�)dJF�uI��ϸ}��E��=�����!w>):/��E*����ņ0��^t>��Ǝ��3^��̗	���&-�P]�K�P�c{ʑ�L�zW��v`����X=k�ʹ�#�h�͝]����ؐ�%Y�$��7(!H�l�z�9gq*��|���_�]����l�^����@Q|����fi-�-0˰�tH%J:�s�_���l0d-��`�Q���AL��1�K^�?#�
3s2:��J�iѣ�����(����������:W/�> !�)�*�����IѨ�O�^��s����{�p\/3c�q��1�Y��84w�.�����Uhd�^0�A����	�<��U�G��~!��������8��-7���3�>K��a�C{��m��aW4VT�e�͒Β�6��7 �`�bmk�A���[�9Y�ҞAM���oH��F�[��J�O�}`�̘��X�f��)���g�l���w��	���h�/<^ǸT��ۛӆ��M���������P�|Hu����ν��anGL6m���ʌ`�E�64?��&-�+U��'x���m��|A�_㵴9�R�}M�]|��ͣڍ}�U�.��!�v���U��&��f�ڼ��3�(���?c���*=h�=)b*�W�yJ(a���p����S/ �Au���ODٟ|��""F,dO�|�j�	)�Ьԡ���B��F�H�U���z�#]����,�j�r%���������w�>���kz8��y�����;@'�UZ.�D���;�큙v[��3�P_�~J�+=}"�9�a�rl�)B<7)�d�ld�X;�J<�t��!}i�	���67'f-�,�\~��e���QY��O���^�{���p"P�S�-�;���H;�jN��������zGR�����;՗&�Y��-�h��]{�<����M�V��v��N�Z�x�y/�v�K�Y�i���FJ���Ë|	�~\���	�<@N���W���D��A��� h��+,:��[��G���YщPf4hOn��b_�}��Z���i (��/[�#������@�=
�G׸/�����Ǝh�P��_��gF?m���Ux��PL��=u�\��A8�<�U�f�#����߼����T���|��u�W>hlJ��sքjn���@�@�%�KM��uc���@��crB4-�S��϶���=i��
Y>\m��mxJ*�kp+m����Y��ikj���R
 �����7�_-�23M��A�{���u1��q�E��<3�R����F:Ѳ\�!Qp9k�p����xR�ۦ?���o��^�4y�u-H^E1��T��_���*��Q|�X��^� �x;_�w���5����ݝ75p��( A�	�zo�$�{ ��qB&u��ח��
v�.ha����J܎�ms���˃ J�aV
�^��Ms뀽
�p��3��a�F�{�8EQC��iVRY���ߥ�1��v ܞ3R!���=$Q�Ԏ��]�s� �W6:�N7��@qQ�J����b�]��Pr5t�RPי�:�'�T��O��L_���]���l�?�v=��7�kM>b�YDb��b�c��R��Xѵ��1U)���^�[b�eE��0�_A�ۀ �0�.��`��U�P�_A��r��w���{��BS��=l{��o���C��A��IB�� Y���-�=\-�3I*��,a#����^������zfD鿠�")�8��5&�����7
B��c�ќ���7mIXd�H�H� �	����t��ʜ݊ULHu`fc��3�e�E"UL�6N��� ݙ���I��1���p��`�n�x˿��퇔ϲ�(�M�~�wCv0�=���!��2��qO�T[$�QW� ��E���vd|$.Gu[L(^�1���-K�j�Y�/���v��������?�W1Ϻ5hL$Y]�����'~Z��t��&\���c�^����j�I�%��"�IhiC��{���]��
�S�y��c�hY�2�,�=
�J���(1VDS������eӠA ����05\��NFc�.�[�w &��(u� ��W�G̷v��G�Ғ��Kb�einԈ�YD��C���ܾ�� �R
�S�}H����=:�7�}C`AY���\#�҂�U4�tp��Y���V����ӸB�Z�v��(lW	+x6x��(��f����Lw�~�ǭ�o`S� �-j^�fsI�)��q�����u�����������7���w�����
�ƥ�iP�,��}8~C��Hs�d��GeA�XE��d��d���o@Ut(@�]������9�2�ϵ;mM�9���m�K�a������>��T4l���!�vQ��Κ�C�7���a1����d���"��,2���N�H2vgmi�tT'�'ܒ0����?J����

�O2�ϧ��;K2��RE��B�6�Kgߊn������QT����+�9۸#����n��!)�uaLh;���c��r0J#�(�&�`@`(%���ʩYB_~��z��
RZ�oE#�6Я�r��uP"r������^\�� �*�ߡG�0��D�yϢ;�qJ?���D�`���{�����s�ъ �x	�.����^+a],<���&O��s�5��oˬ����8���� ��_켋�mת�łG��r����Zu�.��%� SBzak��=ZMw�8�O�y�*:�F���T��,q[�؃��7��o1�6��8�{�# ��(dƛ%�?fza^� ʧGث"ׁ���|�tg�w�|�"3��qE$��F���T.l�v|C� Ȭ��,��nOm�4�]���Ա|i��A��Ŵ��� 5%`�oGg3��Zh���-%Qӻ�ŕ����l�"�1��R��wД���7a�P�=�1���%m���ãT���u�iMy�i�-'���x�Ԍ�!!w�KI,~�$�#j��6�jZe�����ׇǱe��+�P��H�f���z|J�OPsZ~0�z?5<��$h�3د4a6��
��ٔF��?\;#P�)��e�/���=�>I��*��H
ޅ�.x�P��`ȲJ>���M���{��W����8�8�'�IV�����jU ��;d�1� ����ր�r�_�7�k����	�^<,B����3���0�|%���Am�er9�Q����N>e8��-nصR� #w����1�@��+��	b��y�.ËlO�Մ˪��i&;�~�h�����}�Ů��Nn�������#� ~�vۅhj�3\6�S{rA*r�KT�gG|փ��@g�8���w���"ܸ$���ƐM~��q�A��?��%�ŉz��?z՟�p�w[�dDs�t!n��8�*6I�i�3{؄Ij�j�8�a:�:Z����Ϯ��}�z�D�J8��O�t:6����kK���Y{A~����9D����
q���.�@�E��;6w�{�1�㖮�zH3��Z�2�^&��<������%�4�az�*����:	�=f\�F&=�*q�Tpĥ Q�P�ן3��]N�����{q���<�6J�����}��rP-u�e�1$]�0:��<^��