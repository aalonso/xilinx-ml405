XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���f \��M�	�|��O�ρK���S��4��ع�ʈ��Ğ���2[�H%����#<��5���C���J�o	���i��7:���
=��,<���*�Ў�5���0�܉%?"�$�<�(��+�~~'�"���S�,Z9����hG_�3�q���W���:g�>�g����s#�=Q�-�fC�k	q�.q��/|��ff�_�����ݱ�����6#����/Q��s?�|x�����{�r-н�g��_�U��U1#�������B�P?-�Vg�*�UoThȀ��(��#@Av��j��q�UZT-cĬ�J ��O�"�K��:�$��+��\�Oh �>V�/#!�)�Y���?1�pn���a�ƕ�M*� 0i��L�1b�؞��5k�Q5�u�M��u���'��s�	���\�Y��4$��ޡ��Ӵ��m���HOaI�7�
��nk$���/'�z���J!*C)q���N4H�\(�z �r���v���/Q���ctY-����I=�u�7+��'��ѥ�Q��vbc��/�B��AA�W���lI���9�@�������!wM6W���;�������U��8}����=CM�T:D.k�A��8�?��g<^����^��n�_��b��\<����1�>;�2��I�h\�~�{i��3�3M�[��[Ji��DWu2��n��M�[j_��i̋��ο�eMW�rL���\v�ER�\J��y�v_@H|��Z�XlxVHYEB    118c     6d0���L��O7a���F
;T4L `��nI,�b�W'�4��݁���bQ�&�P�vQ,��K�Z;���H��=F�}c�T�LjBvߜw�n�sM,=m?��W�ߡ�r����/�����M�Ȃ�1� �>��F���C�~o�z/ɋ�������f�1�gˋR��]k��WD��uFaY9�n�������;(�Qj��G�/��D$;wo�Y�u?$���N��` �ö;��˾��y����Z��Z��	��a�*t�'	h�����}�^`�F��%�6hz0e	]���؛����O��\�%�{5ۉEj����p�r����LYw��Sr⺘��r�˜T�'ޚ�+�_n���&��ҫ�<\����Oxú)��D4��i����J̈́K�:�T���Lp���*M��٣S�ݴ��|*�w�sd��਺\k���}W�������3�4� �葆,�f"�y��
�+M�|�)�`�ɧU �T�pL�/%Zxj��2'C&l��m/��w�J/��xB��Wk𘔎�{�(���-���4�������F��fOޤH�Io��{��j��b*3mb[q��8H7	oV7?����꧊�����(�W��/%��:�U82J,0�L*���U"�eh�"��ԯ�Y?��)�4����xᯄ���v7���֪ťt��5� T��D뼝��sJS�}|+���qٲ�$��.���5�C'5�5{�P��X�4@wJZ���=�*PӴ�4d�3��{�-̓ѣ�(��<�x�|#nu��	�v�����4��~ Y�H0m3	[]�^s�^eF�����ʵї#GwcI�4)��t�U*��r6Ak4+_��G��c�Z���z����	��Ss����,�km�����%��p��L��*X�C�A�s~ӈ5}�}��AjS��{>��Ò}����a����eS�V��j��s+銅�U��?������l���p��z�jF ������C�y��F���
)L��Jϳ�)�����X�X#$�*bQ�&�}�:����=�������j�N?���[�U�2�<�'���p�?̝D���k��W:�]��s��\�r�ѵ����u3�K,���3��%��,g��.!QAGY?9
�LM�B��j^�Tڽ���0�!n ��{=�b"��f:�E���=D7�IB#��]��>�cz���;DO��Pd��~��i�b������Z�����l�И9�a�`���T�u�OkP�ԯA(k��Ɯ�3k	�W[���+h����7����4�%+)�m�D`&ڐcG��*�Ii�Ѱ\Qjn�̿1��Qc������eQ�h�޺��ۃS�]68��{��#Q�Y����.wb�t���"����BBhd��X����K
����sj�XՌ�Tl�?��g������ϵ*����Dtc
xC���$9�󰰉=Eh<:c
aV2b���Ƴ��mKQD�A�'�eٱ�HrK��hc��בG�<,�¼>�PF���0Dp~icr���ş��^ <J"��J��j/s�T�BJҬ���K�<�f{�E��I���+�tр���X�qPK;��;O���u�$�`6��ȇ�?�a.�X�����qG!щ�/D.f)Q��\�hʢ�Y>�s�0R�k;����:��IeC}R����Ah>	�����y�>���	))��	�����	�{{�A�>���E����+�