XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �<ܸq�l��Fy �F03|ۑ�Z��I�T�ҕI(EwR�$_o��P�\�QA�r�I\c�8����'4Yb��?ɤ[���U��6���៕jվs�L���a#eM��A@����xhR�
�tJ	����T����������],��9>�V��i�O\�WP���vU�s�xk�?��׏u7G��vFH�m?}'����LW�E���2��I����D��7�4z�~��w� �d���r�>(�M��K*Щ�6��~O񧿋ex�[q(����8�T�y�Hn3c	�i�#��3{c嶩���'�ޥ7��ш:"�(VE{�N��&d���~��J/�ɘ�t-@���V
ꗭ �� ���|S2��P�oK�Y, ܈�T��6�����K]{N����e��෕��M6FP?lq^��#�s,�V�=����2�Gc���-�h�d��!˿'��G/�J��KC�l��y7�ޔ��k8����D�{Ǉֹbf����;Ee�j��7Hw��li�x'�h�2la	�1{ջ�X?���2U�mW��U���A��z���b����X�p�ſ���f~�-�&�^(��j�˽ު۩G��2�n��8`���H,��
�Ea��YqP�t���͌��sT�T�Fq�|�A����jg�D��v�tȈ~���M���6���m��T:�M�N��iXB��Xr���j��+�h2z4��<?R?�R)�j�ֹO��z���h�Ml'�@��Q�x<XlxVHYEB    3f19     db0�a������+��_��J1cz��I7q��p�I#���c�����Wu�Jk�9:��%���h�&�`��$���βd�M�;h�%��f���=`��pG@��ob�/ �wZ������o�Le$�u�@F�yɰr��Ӗ'�)!+9���Z��o�M��҂Ƅ�8�R!F�{d�ܓ�ċ���ԃ�èL]PXG���@(o��{�{i�����=�6���i���җ��*�{���8��^�=�r�_�s�^GY�V��9�.��3a�1p$� ^�M�U�B��W�Ŋ�Q�i"�$N�l�t�+֓?�*�\S��%H�X�6�ؔ.t�w��J����9�&rG��$Xh�o��t�<M���m���y�#Jyp���;1���-b�%Q��@^^�3/���U$=t)&�b�H��ae�����p[ֵ>�SʙOx�K��D8�I<��^��f���X�8�A�+ږ7�v�������$��֢ O�3{���aD놠���&X��0�
�h��n��������І���,�1��w��Rѭ��q�2m�r�t���@ްg�~ ��6�L�y=N5�H��^���Vл�z#�F.��a�"a�Nq%:V�1Z@J�y�DO{k�S����J��;�K�����Ur1�e���cs!���o�I𚽜L(؆���������q0>'�GQ�"��=�7*@��w���5���a,�}�} ��Ր�~�x7:�Cn��
����<Tk�r�ԤR����c:C����3�ܪ�ˉ�f-��5z�i�h� Wv	V����}|vt���y9Az��4�(3j��{�#�~'#g-9���Mw(�?n}��/��s�b���X;a��
e�Ӏ�1_���I��� �n�"��%sS��ʲ֙��6Ȗ�?����Vp[���4K%��Nd ����oz�xF�M����eٶ��i+����UV��>�d��df�p'x���G._)ŘU�������>��A���T�Ţ��x�/�~Q)zP}㕋*��#��t�<m+��?/;���o�����:���A\�k�p�D|.Qz�M�d:zx��M����ǝ�xu�G�^܋���w�gSS�R���7�UI�1v�+U3QZ�Z�25��+��&֎��չ�:jDq�8�[ٺ�E�U�Q����ށ�?l�y]�Bx��}��Zl]�;2��pl�v�~�DvAC�8�הoh�ִ�"�Ʋ�7�B���qHW ������
�U��!�!�Y'���tl��X�n!���H�d�� �~�t��W`ݠ&��Qk��LY���r}�LG*�Z�>ȹ�'Y^,����3ْ~,��	������a����`t���4t����GT'<T ����(J�AUuVë]Iy'���Ԥ��^0�c��V��9X�����qg���T���(�PfUY}�M�������8��#�+��g?Y���)�py�_��Ho~0�����.7�rJ�}�^bW�d>[��ld��]���A�s�J�˗]�ۏQau���h��TK_7]z?��T�K�PJT��n&�&c'�y���y�=J��-�/B�^�0`���1֎Nˆ\�I�8(:�����З��׵Q�'i���l����DPeB��㿄{�e��8���ԂpTt�H6��f%�(lNtg�v,6���١�A��X��~ß+m���1�nb�5V���,���ʻ�.��o����#<�##��%��G�Kƻ�E�;PF�fF�ĸF�
���e#��m�P�Qx���7��+�3Dx�b��Ĥ,RUBg�~ ��}�H$���(>6�o鎇��E�h%mj�RB1;,�Pp �ٶ$��E���Nǿ�i����]�py��rB/�k�N�ĉ��Co����y4�s�ib-�I08� ��G������a3,@F?�c�X�n���Z��oBaU�"~0�=Ha� �i���y�u��M>�Қ�qsR%P���sNW��燰h�R������cQ0J#14��į(����l�_��xʢ`�J��2M���4�� �f�K�|��C���is^rE���7��r>���0Ek�-��6�%� ��R�xav�R-0���'d�2�&��a����RSYo	�zE*xnW٠Ϡv�lX4Sa���t��p�Xtΐ55��7�BW ��[����n*FC4�aiy3��t,0IM����:R��X�G<��H�B�w�J��v��-�A.����q�4ue{�����h
���gt��&�ۘ9Q!�s���x�����C��qT���|H�+�3?a���u��'�7-u,C+�(8"�ѡ��дj���޸t�0�7����+�� }�	�{L���◶�G*QEj�G�����_$��H��&��c�/�l�+8c��垟�do�s�����_��^ݐ9-��Q� ,�F�k�w�� ^��oIAR��x�bQ�U�B���,���V�e����S���#<p�E��ה����lq5{����5��V�n�{*��	��UM{������(��Z,�EP�k���1Ȕ^\?pp�
���1��\V��U�K����{<��$>�ʰ�����.�Ă[�m��|���e0�Gk9�'��Rs��مY���YcW��>{&8oV�W�]R�Y�5�\���S�1UO�+kl�ˍxh��7*��Ed/M�ǌ�0��^�8����۴�* VlR��
�
D�0�U��mFu��ou|�2=m1�i F�s! 3,O�$ ���+e��,R)HmE�E5�����Iܮvd���F�Z��x@�;�m/Iw-��TDb}Z���M���\M.�������r�5N)ʔDU��+�r�X������Y~P@�pfZ=�����
��qč������ �+�_��v8�ɶ�`3;<��G�ē���{���-K3�P�(|3hLw���>�x��)N�ziҗ8����J��Z��i���Zɔ̅���F�Q�&-f,$�̓Gn�LP�{O������l�X;՝<kMo��ȶ�h暈��Nj,��YE�X�~�;�)���C"�]){�$0��In����ߦ O������N�]	���a�#@�����/�> ��(��.�BLGn2��Ck\����=�(Xv�Y,}��-Do�l*�C�e�eJM�5�CS.�ȋ�l����&mR6*�7�}hƻ:i��'�����:׬Ɂ���~����R34�Awc�h+�cR�����h���$���%#�F�����Mp��Q>%ݲ������U�{n?<��e��ǭ�o�
ԳC��s��PM'c����dĝ=�
��W!��!өJ��^~�]���r���� �3_P��p3!ŋ��-��t! * GT%q���J�F��Tݫ3QMO/�ځy�
��9u@�&��[�����a�9Z2�\I���7�a!��