XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ѯS+!�c�s�W�FM��[�s��'y>��ia��J��֨8��Uw}������>4zB�>��4W������N����2Y�fW\Cׁ.��~���8�H"���'�;���9�8���o	>�j��� �H��X�;=D��d�d�ٺ�߭�uaJ��Oޫ1�Yϥ���x�?a*s�_<�s�Gֱ�1��ΰiA;@�mDV��*Y�����\�YT�B��Ѭ5�����t�.�����|:��k�оQD��p�,B}QB]"O>4�(���pnq��#U��9	��Ɂ!����Cɺ~>q�hw��%xe�[�!�l�>���y!������R��}#��1(X�-Ui�>B��"Hiy���Mm��x_�II��G�'Cԥ@g;�����$�WcV��V�w]����=�j��c�E�M�)_��Z2�]z-�\�I[GQ����Ճ8�3����W�Z]lv���Bn���Gs�.�>�r���آrܒ� 9��[?�O�*h�%n���8yr�<��F�2JL�`�)�7�V0}��^Oa�%���29�;��'��FCt%y=�~�����'���]��}C��`k�t����*/���R�*rg��ɧ��u��CL����=[!$�>lxIq���8�tP�����ιWB�?�&-�!��W~��*�X>nAoے�F��L�yR��Ĥ*�?���Z*-m�+��#��/��ϋ��h�ee}$�a��~�-�!��#c.ڤ�ě:h��L� �����7�uXlxVHYEB    4564    1270�-�
گy^,��ghd�3�)f�PaE ����H��,�5É<S*��o���2��{o�Mߨ�
�u���ջ/�%8��F�#g��l�1�03H�������݋�D${n�_�X+U��3W�=�s5bz�/����U�)-r��?G~�U�o������U�����ˀ����M��Iot1�xi�_�rC��z�juu���4AAD�����;3�� є�C�Hcm��F�zM��z-�bJ�
�e�4�+�01b������v�|@���dk�e)�?�2�t#�Tz�1Ի1��?�UR��ٮ�����7�x+{�e����������#���BR��=[�yՕ�]a:0�:V��1��o�%ɿ�����ag�{�[r��'���^P5z_�SLHwC��8��X���V�m��D��Ue����:�5z���I�m@J ��+k>
cz��:c�꾩�Y��b�Z���,`�u�CB=;F��gM�R�0�� �s�OcAB��V#�M����xOk�0�r��}n�к���$Q_9�'s�����f�� @�p���Zg�`O�8e���=�/�VʸF6�{�G�ZJ�0N�f����l𱪠���Wu"yO��7�E�	�4�ڷ�t�;��xS1�k:���Zw&g�b�����LN�^��ɤI������"2L�^��֠1�HF�H�Anyx����.�uƂ @����&�P�+%�|]�Y	@�R�`>D���������	�4�
'�[P�1^���p�iM+埪��`����C�w�Ѡ+�"��ߛ'>z��::
��Je{�:e�i�R&?\�O�R&K���6�&l��k�?�	��[�-p�II�pa4_��1�
�P�s�#u�m�c�h�M`���;�H�X��!V�RU��Zg�}m����Ꮓ"�M�
�<�eO� �������7uTB@�1|�%g(����%�����lz�&��#xn�ԙK���$�B�_�t��Gk�?<�&T��W�5��D�!E��lR_d�I��(�|�O��.�jj�S�ߔT���U0n�B�DZڌ��U�0S���[o��a��y��K��O?A��5�O�3�Õ��aW�z��.�UNIϻY�'0��|��V.o���郊�¯���a3"����͞��k��U�c�e��:-��RQ�֎���\8��W{b͸hxܼ�b�m=zzi/Wy������1�;#9����em�I���������$?\,��gC6P���p�.��C{� (���oX�F�n�����lN�KHɈ��uz�؀�8�A��k\�	����7�%�D�g��ڧ����V6Haǅ�m;��`�[�}x"��D�*Vb;�^�x/����D��#�%�$�� ���ʐ�"7��׽^�]����ϑ	GZ (<~�ܫq�[�.�a^���8쨖��Rw�*K�ƥ�*�D���V_|��� EX���N�0HѴ$☾��Y�B�x m9&/�)JW<�R�e;���b�����B'7wu�>���!����}��xq�V�t�3�gZ9A@^�%{u�x]$�<B�F@ 	�%*F�km���3GN�D�� �b�؜J��u�^KWH�cأ�ioe��<�W{��i��)S�F����5dw���ͻUT+���1V���������@LmR��|G�r�d�l�H{ۆU[MENo߫����S1
�ڸ�p���ّ�#��nȖA�������ϓ�ir��g�L�;��<US@�7�zճ���;nE������,�a� ���w��2�^:&����/֋g,�+��>%��?P�W1��Q�6N�AP rh3�/���1]�
)�A&*m��mj��F��)b=A�q!Px�~w�rK��P��l�ۿ>lr���=��3Jk ��6Yex���:ܼ]���o�i�JR_�<���|��)�>�x/����,�I�"�e#�=����	��m�U�h?�����Z����qs�Oԡ;<���dc<d#����3H3�㧡��#>��A�u�,p.�H�6���w���)�ju��قa?6��v����~s �.3�Q$|"&,�����ָ/�3�lFJS%Q��g�E*�8|�I򟔅���m��E]�����}WÞ�� JgcG��#�Ї%H��U�fCd��@����
�:�o�Я|����͇p��\3t�4�6/��$���B�\��` 흶�`�T�Ҍ��?�g���]����@���..x:� �ͭ�U�k��ȶ���r�j��w�S\��e�M��a�4H4��*|���Dv~���]�o$��id�kr���������2�����ЧKL�QFid�"h�� ت�ty~2���B�z�T���K:S=�#��Ç�{!!Vo8XR4�c���K�fIζ,�(g9���i _��7��?���\{�v$Q����w�>��r�ű⌔|<D "z��O��t]tۦ@��̼7*�jH�u��\��1r+f	8c�����=F����Ɉ�?�of�#d>�[�[L��TGf���7OW�t}7����u�i��1��O1��1i!Jx���ڸ�@,/�i7o{7�kҒӉ�-X~��(�
�r<�u�	t����hml�\��J۫$���ȜE�FC�>IZ�?pqHT}	��e�xO����Sf`v!Y7��38��y��j��H^���O��"�Q%��%�8�g��;CS]���?:a�if|����7�G�ĕ��H���y������ê��!r�����Ѩ�Њ����x�M\�B]/�y�&	`jԕ�'����G�=/9Q-X��bi��C[��9�Q�3k�G��] ��@�!7>Q[��<r$f{�<�2���d^�� b��1��3�$�n����1��b^��P%O!���� ��{�~ռ9�3QMuɼGȟk��U�1M��c��p�"u�<��}���9ém�!?g	�W�IiY��{���;��N��Q`	j�l�]�) �f�[��
�b���O���yP��F^]����<����K�Jb�p3�u+ .���]�J�B�T�2L_�,�'W�ul�8{����J������uJΥ� ޡ���J{>':Zp���iLY�]̒/.!n�i����W����8��v�A�,M�}$s��?��a;]�A��������"E�vq7ߛ[�\�}pH����"�i��ѵd��;oC�����>)���I�K�qکX*����)G���v��*=)�sm�4M:�I>k����I+�2��CDY����^�k��8��f[z������"Xτ�)3`���`+EOLMr�N,o�F\�PI����9c���p|ԍ��F2r#�(A @<�Ǉ���l�{"��ᖻ���v�E����aZgI�3�O�:H촾P0�
�'�M��+�%�#�:|>�4P�lwG�=�أ��yb�}�f�:yƀ����6,���;נ\������mt@���[E�P��o����^���!��� ���-}D��L+^8�V��ݡe*�v�����
W�]*z��J��4�g���y��ݑԶY 2,{0�.��=��eO�j#��� ��c���>����2�?�A���+��B0w`�Y���r'��n��J:��u@�̆ja_4��D�H��'D
���i�]c�nN��W.��T�>��AWD�R.^u	F�5*���:�`n�����Bt��-\WET��#+z̯a]��=ln+k>
󍤗����_� tJD��7|�T�uI &�m�fҾ=�nZn������_��C��e��p�Fϰ�b8?@�U�;�t�YT�yl�GJ}ڤ���z�@�k9�-Z��6/�0j;��_IJR.���K{�c���INnc�w���!��o?���;[q���$�&���c�棩&��)R9���"����6b�o�~,�O
�p.�"aRT<'�44ފ5���Wfh�9�:���_MT�5�q[�D�y��3(HH'�s�rI�a��_��ۀ�y:p+�xM�3)0ፘ�Hh�������P�m3]��A�9J�@b��=�~���%�����=ۘm����N�b�����7^1�u#�8�7�u�BF8���@��{���r��}'jܴ����:������a���>�(��)���c�����_���ҙi�.�rC��d�C��L%`W-�ľb���j����\omꎏ��|^��Yݯf�y�i&�I�j�F�Z��M�6���Z��0s�[�2�Èps��J���yM��mAr�H��MՂ�4�c�-�y��)K��H�-�שn��=��*�Hm0hz{,Lk����I�Ê��CǴ�+i�I�M����C�R��U��8KSD)�z���}�:�{���t��U���%`�R��q���G`�O� ��&t-�ppQ�QE|�b֎Iۥ�9�M��7�~?!�C��r�K�'��0.��}�y"���~��Hs�-����ϼ�+Vk��.,Nc�I�+��-�V���˂�����~��yW��C]���+�;��_�9I4��y:9�i��2���tJ�BɅ�z]F>���L�2Rl�M�v����Nހl�װE���|p{w�и�`����"j���ù��:�����%��H��h�?4�5�`�����B��+�yϵ���*����=C�cnDq�J���Z����N