XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��mD���y��fђd�|�ζ�$v��	�@w��q9�ו��[u<�B���D{% ���k����/l�e]�PL��]b��1 �p�W�J�^E��HMW��W$\����+��>}�I�e�rq��θLSu{vyRPd�u��O����I����_�R��!z�v�6�����N�o�؁ǿ�#�Q�9�v��.L_����09�/��ľ:'��u�,��BB��n�͠n5r�=�7J=V��XO� �\�����]x�_���LIT���,l�!.�;���Z��)�l�8.˸�!UB_;���(�wH-9-ڐdP<gF0��ϞCT�kM�o�p��I2�:2�O=�y���2
U�~h��C3��_�E�3���B����fO.�1��wtK�
�5;��w��p�a��r��'�m��w{�.�=��`�ns<?B�A\�s.��lͿ�y��`ۭ��8B8�Zs�'&��=f���1F��~h!�X��$�K���-w�̴��,��&b)���آ4�1�b�K�퓈Iً��TI��Hq���tL�$��d�~,��hH:�E�3q���Ԭx\kV"H�c�Y�q�vhU����x���-�g���A���B�@=@{,o?)����&�6b�Bߡ�u��d�X�<����l�"�)�
)�Z��M��b�f:J)�*��`.��Q��Ɛ�z�å��b�{�@�m3�
h�B=-5��~Mq�@L@/�%Ր�[�?�E�~T�lB;�B��R�GJm�XlxVHYEB    6ff5    1760��Ћ"�aT�6���� h��S�ǅ�,�V<'S#�����	��ó��#/J6	K�Yץj������Ɛ �-z��!�6*W�a�! ��8����Њ��Ƒ��xQ~��%l�[�D�O>�Bk^�aV���͵�&��Z	 g4����臓FTJR�KćW�y��nDՠ4ֶu[tS��Pp�{@��x���؅�h̥皟���j�3n������#_簧�c��O�LAp���n@ނ �]GJ�S��%�N��J!2����3��r5�$A:A����QJp+��dj�y��Me{֍�}`�@?��Lhk/ȸ?ɐ��� ����[խ��Q;G��U�����k��^�� ���Y����˓�����P����	�$��5���Z��y����KI��R�U��1��IO�_�G}[��3근���\��D��7�����{���	���Q�:�����g!Y�	<�n�p�z��� {��AP:�F�ҲK�V��r��;	����.�L���ա�����E���_+*X�����r��Q=�c7wXJ�����Ob�G� bH��dsu�B0K+�/��0"KIP��@�@.�"Gn���x?�f������'~f'�"���T4���"*��7�Y*��m�c���}����.d��,O��$��q���~I<U�>��w\���8/g��<f&B���!��:�@>�s&T\��RM�Z��ƗG�mPl�L�B�{�b���J.���L�1c�{Y��x�e�q21J��<�q��{7֣8�V�@u�9'�ځh��"���B�2���#e�y|��D��RiT<37����k�U�O��:.s^�Lb5�}��	�(��M���:�Gv%u*�j'�����3褠�{������N�qj=}��MI"g\���X�dFDb5C�35��Ւ�Uv��q�{k���gg&/���|��X����T�@��7��w��Л�-��6r_� ���{�e2}ۀ ��]T�:�ʷ%jib*��W���9�����4������-�.�/�����l��7�s�T��F���\���x;�J�ՙ͊���S�*s�F��+�x�"��?�`�@�&���+�:��.�4D��Q��ڶ��D���#�<S��\)�U�WTғ���=3�&�ו�j�}�ŀ�P��3��Ye�~���>ُ���ָK|�:}j��M-����貮�^���F9���/R*�(�=�=���,��K�t��?a���`�����"���B��r�[�0h�����<��AaTFl���������[HY���F�p�Kd�W�-6���B�q8
�N�}��(�/�c�����]���_L݁Eap}eN�h�IY�a��|��d\TV���.�pV6T�P b���3���I�W�ڐ>I���$��?�D�_gvE�M�D����`�Ɍ����_�vH�C+��H�8�]�V��?E^�n�\2�����KQ���㙟���ˬ'3�GD0�
߶&j)2���5�*_�����O[~��?��.V�T�HЌ���Ъ�Q<��Z���(Zظh�&`f��~Y7;�_�B�o;��Xh%W�$�=e��穻�ć�P5!��KN7WmEh�i4ss�Dlo3�1���q,oW�Z죯�i��.�4��7͵��C�p]�I{2g�iG"������4��w�3�CS�⯱26���|�:�����WHA@�{�/O���s<t|�dt��r������8�QN����j�)�?�Nꏧ�	����?�9�Sh%��aK�1g�	��Ԝg�٬��1��&�i��J��7r΂q�^�Z;���#�" _��><xQJ:P����ѱ.\9	�XP�<�ɿ������%#rNڳ�7�����/���1w����g1�#�@�����*��Ҏ&(���sKV=�A��R�I\��r��XT�}X�u�ß�T�|�W�:�H�n.Wj�~�i��I�3O<`�le����<&9g�y ����3/��L�6Ee�3���+��w���|g�q��N�yH#	s/�6�m6ő��/��+�
�;��(�!n��j������1y�$������S����҂&�T0�M7�4}�I�POR��%n%&]�Ư��q��e�H�E�qY���uQU���;;�6S��s��΃sX����V��c����9��rlI�&c�}�H��Ex�){a5����';>|�V%�z��;Ocj5xe3
� #$��o�ǀp�?]�����;PF�� �T��uȒ�jgzZHWK�-շk�~7�y�脨"���-��*O�c�ua]N�9B3Q1����:�r��%��'��2�|��%���5nԒB�X@zV�.�9Šӝ�ߜ�{��,q@�g�	eb,�����?��1e=	���1Ѕ���V�R7�6��°w�l��w"�j��^]|=<�����@��P끴��m~t���C2D����14C����T+<L3pU���pkQ�Â���`z.�1_�t�H��%�aρzB�I��d�b+	��Yt��0�&V7�U���lw�C�q����k����n%��K��${�Z��oc�|���n�QӯM� {�9�B��$~��t���'C�W��v�l,�X�<K��]�p����q�*x�m�
��вh'�p�d�{��pN�:�|�XE�+�^^jb
U��!�k�v	��uW���g���.�0��p���-�Z&nE֯d(�c�<Gtse2�w��Yb�z���K�).ɕ�c����-d��\͜�qEo1
���߅�(�8G�쒨��6��AǴ��$���5��*!ﺳ�g�����6�P�f�]`�J5?# L�Tԩ�ߍdӮ���8]*�'M��'=�f�M�yv�R�~/���Qr���)I�g��$H�b�_��|1�	5W�w�+�{?�K$�`ś���y§(�*@|���03J"������U�-�C��+W�w-$U�n5zo"��;҈�TM��9Q����y=��R6Ss3��Qb��L`�DN
 �7v���a Y�<S�%�BQ�{�#���uD4�_���e�.�48]')j�ҹ�s�1�!/G2����e~�I1j�៝x�+�3C�V�aK۹���>�T�jv!��L{�{:�P�4c�=����VXV@�ĮeIx�m�����q��_���~�)[�g�[*J��x5q�N�C��<dY�T�igI�J��J��P�7U��?���跜��@_�sM<��Cd�mӅ�[s2�֫Z5��T�nd��Wx� !��I��݉Ҿ�5�0�'�k�)UMX~E���HP��K醴f�9��vzS�e��xE-�|q]�#v��3,�X��Q#!��N������ȸ���Zr�����%v1p3b��q(7���,'eK�uN���y�.��y)����	��z�{-IW���0��H+�hb��u��z�����;��32(
ڄ��W�O�e��CkkQ:��I��r
�C3���1I�@�����B7��Hh�ǻ=�$�+6�����$;�g�}ҳ��C�֬D��{�ы%������.*�Z�3�YC��U	�����9tp�`u��	3*����u���͘�
C1��*hC��+�L�*�!cT��mt/��%Iu��`�G�9A4���WCC�5�ڧ'O.�ȷ>Z�b"��St���P��]�����n��Hnյ2M��������Z�	��Hݠ�?Nl�
O��|{��R$�f��]��E���c�?��X��սc�g���	����N�V�V1��j���I@iS�}z�*��c)�Y���i���\Z��|ğ�)�F���ZG�|:����̒��{����P��T�U�Op<]͊}&*��Nm	w�����#��:�͋����.�ǉpj���YKl��G��Z�!0"	�/q>gz�Q��+ ��˶U�{Q��\0��>eG�W����iw�-7�|�h�p-.7�{�r�����{9��;σ� զ���Uƺ�8oǫP��Q�x����|�@��&�"�h�{w_o�Ǳ*�+Ms̞wV�1���A�XS����2��K��z!�γ\c�w�!A��z�&=�"F}?�y���-�Q�A���\X1�T���Zn�!�Y���K��#�b/��b���,�/��n3q���(�hF/��e��.��g��&�����V�� �̕j�7a��7 n w�T"�c^O��P75�ȓ7��5^9S��o�� �R��l4��za��&��3�O1C���ͣZU/V�Π {~�H_��F� M�|l�{�Ċ��)̤>�Q�v��}o�v�nVnwr���K�:s�J�����1������*���+�O"��:`�?^�w������)t�`g%�X[����;�x�ӽ���P0Is��ݎ��z>/i(RJ�-Rw�:�<��b ��A��bc���@��S��o����4��%aP��vH����g��lgL�	�ٺ�a۴xdө��yx��%4�F�x}��IGU�i�j�2�g�QJ�U&{KUIƟt'|����6��$�Q��W&L^��]��d���.� �6�:>>�W�f�0��g�����L]��	 z�<F��r��]�!���գ�7Es�D 8���/��6=�I �wq{�EĮEZB��eg&K�,������Ā���&���\�'�*��������O9o���M�4�V��J��[20����X��|�K�x�I�Ì.����(ٟn�F\G(r��i�+�u*%�uR�N��Y�`��W̒��(Iҋ6�$�eZA��he�[����,:������_�,a������C@�@Y1���ˉ�e��lK\�`�˥m���}���Q��:��7�紿()�ذ�Z�(���ef��fX}  �dIɾ�ka���XHXTG��7�g�Lr������@52)[���G<��p�'��~\�`��~�R��$���u���C�oý�I5��e,��{���E���)�y���A�&8�[��R�n�4d��;C���R�jf~��!B��y�-j�pM�3E�4`�+�M���3��
�7�8.�C���>��\��i�fS.	9M�^�kV�n.��i�{�k3�� 3�Z�2r�9l�6$J���-E���tR6D�ڟ�ORm�̲!��)$Fd&wMY���Bo��0m}!Ȁ�{9�Ի�@��""ʞd��ي@1#f����������=U���;'���� O�,Tt%O����7���Kb�z�,+���V&��1�!|]ߩPu+I�59=�⿅�&�RyB�D#4�j��L!s�q��F���C�x%r�
0z@"��<�㢮�XI���6[�щ�OS��`�c��Ə����gI��N���Xb�7�k'�|�
=�(3Fg M����Y·j4f�+A"�6T�'�����M�)��@��O�adY��"zȽ{��Һ�����4��������e7<�v�g�� xPZ�\��m��C��k���� ��������iB�u�y��8��A�AJsv2���#�݀#v���%Ŗ �=��un�G1M�ߺ�z�����.:���J��a^)�:X�wV���	�t�;f�N}�����KN�j��4�x )\�Ʌá\"OA���}	�d�{�Ȣ~XR����V�)B�s�C��k�ҵ<�-O)��ot��Id�P_�'O-��R@ll�c/�
��0�ގ��{B 7�g\j�9��%�c���� ����)d���D.��TJ/H��Ǯ��������ê#������OK�۰��ol|�704�G�'��%���?��_����kf�Ҵ�v�����n�J��^���8<�v*�O�]