XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���K���Z��%y;�k8���+�0���3�@�P�R�Ch�+���t�f�(4��pO�$đ�Z���y�	���
d�X+A���@�<���(J�1ձ��C�6�s:�,�¡w���?�)	N!��;��U}��&n}D�[� �a�&���xsh���R��[a�[4��2d���F�߻RDhL���FY�]����i�9c�^��q��|ő�D�tY��m������cϷ9��ue�wp�"t������3c]y
��?AkB1���iNW�/?b�g?��|첿��}饪OK&�ԭu����Lu�j�l8���k�T�n7�p;Ta��M�}�k�D��#i��^������a��#b�S�횅�wŘT�C(v~���&���w^٬�D@��=�S١1n�:��qA5��	�y�M�7\}$8jܟ�FpHɂAn��w����T�2�� �Ugr$�T=���wb��gL���!�JJ��x�b��I��("R顎�O�z�!��Y������)�%���-U�k;ߍ�vl&:�<�{���ؓEcm�N �e����0:Q:V�:|���:�"o�3&!�1�ڷ M�"��op�cǎE	�hH!�{Ν+��u����>�k����O�b >Z�4�P��?�P�����i�h�$v��K.��L�(ڴk�l����Ǐ�I�a�m����F��$@?ɢ���6zm-�p�M%�����+�[�[�ǉ���u�Ƚ��ڱ;����C�%� ����B�XlxVHYEB    a19b    1f80�N���&e~�|��T��V�{s���==e�@����!��t���o�x���}��b-I8���MR�CI�)�cǄ*������%L�"&W7���\On,X�ZW����شZ\^��^O$񛠳!��������5�x�`��"f�jZR�����yl��}[���� s	��<싟�	b�A�ta�b춐A�Wj�R��i��1�]����4L�ޒs�^����#V���jyI�} V�����1E��r�XQL�A��{�V��v|�`U�.�@���--��ĔN��{m�N`���(ƁO���� ����5	y������3�� k�%��W�xn7�q���q��d�k%�>)��#s����R0��_��w-�ਏ�?��i\�^�������H8�˪j��79"�<�������ٸ��4|=�>k�#���n�RG�Ť�%�p.�����%�[��m���(�/ΏAc�E/�)!�Nq{"�ޓGFI��r���Lf�s�W�"wؼ���'���ıǽ�*����
UΔH$�r��}�t�Z����������������׀�\ZX\��hw#�zU֙��4�����$�D�J�����5��Xžk(M��H%�x�6��G��ﮕ���I��t��H�C������ßu�tԲ�n,��X�-�V5��wS6����J��hU&7�hX_��0���ǥ~Ů�j��v�J�@5H�%eV�Q8X���"��0���J�s����lL�B�|37[r��;t?��^g�����2.˼����N�X;�m2O��o|d �,�4�=��1������9�{�{���B�$��o�rt�f���ɀ���1�q�������-#�s�ᚼQ���ɼ	.��+�oNn�2�#���U:��(��YN�|O,¹�MoC7�^@�Ax#��YJ:@� ���$k���gR�qZ��-e=l
M��>k��;�>��6���2��7v@���]�!$X����G菈x[s�ׁC�8�����ư9cQ����Dܜ��d�ɠ�Y:���0��N�93+����ęd�Q;�g�m�U$V)�S�Ц �� )A�՚*��|��1b�t�H�t����q��Z�7\�~Q\wz
X����/�bD���,V��e��J�k�o�hu� ~�Li���K�,�͠ቅ��1����EF�d��K�&�M�j}��L��<�����K��3�/�7��|#C�k�è�]�9��ϼT�/��D���sf��F�ǘj�&��A���\�{�vN�����o]���j����pI��7�]Y����R�ؤ�3���G��g�_��y��`�6� DQM�z��<�xUχ���u�Q������h7p�n��b��R�WH?)��#������Ȃ��N�5F��-�pw4�&�)��Y�ÿ�q��d	¥���~�N�8�ҩ���"�p���1!�p�D�bG(hh��I*�ڀ��RF0n�g��3��_G�ɦ�X�hM���[t������C>��&0�^��YR]~����q᫺c!�/�#�v�����5�|?��JHk$�#6!��\��R/�t��%����6�$�K]F�'�����2���p�Y�4.ذ�oAr�H��������A+N��HS��G��{c���o�ْ45GRB���6�C�.=!m�=��P���27���g��g����d}褈M��l�� ~w�r�-��J+���&%�@��@[�j���%"sDV�'kQ������b_1�\�ﭯ6y{7#4Pk��!
~4�;eZ1"�>���kN8?ƒͫI�qwvm�?y��4�a
��,�,�+F&Y��kgi *$E�ij��j$Hn��Ҁ�;uų�ξp��pD�vLP)9�]��EP6����ߤ�3�ɵ��0����1�G��`�m��g2�	���h�\��N�șI�ma*AӫO������W��Ӵi��n��p�������e�D�L��.�#� ˢ�4gF�9�t��}	���(5\:�NܢٱbJ_�� `D�4d�k��j��
6x��Ga=fhD��4��4�[��C�t/���F�c�j��2F�q�b������ ,��GKu|�R�GE���ro�,���Z/��m���w��":�OV�y�͸��W�&��i���A�8t�F�_�N��B�JPj���U�`���eJ����97x�+ �q?�/����yAj���N�M�r�Z��f����O3�i�I��;�EW����-˴BU�;� AB	^I�h��PDF��� ��5:�E�ح&�1,����ٝ�+����a�tס*5g�hX��W:�
L���H�X����_���^%Ko�C�P(u���{�{  3!����<�evn�8$������Җ�sb�j����m������1��7U-�l_i9pv�|�{�Yf�:��#|C��6��S�GPr�n
���XW\d&Y:p~;��-�x��(���윮��f3��w���� Z��7X+?�XfM�b��/϶�T�fE��{�1����`+�E��֏��r5ad1;? lK�Q��U����p7�2w�5%R�w���Op��$@Fg|Lۛ֨�,�v�{ẙ)��Ā����s���\�/v���O���mN�/@�MFo ��ߒH��I;PnS)2�=�
����ZȈ��>̷�_���`�9���}�R%?��F�=�N4��������"q&����d�2O6�>G���ժ�q5�Ck=c�u�[�6Z�&�[!m�㈧NI�bы3�}Bz�5��+���޹]��$��W`�(zL��:��\EȀ@y��L$�C��a����(�wc%N��j^�?���l/Z��}�{;6���}$��D���e��c�l�U���C�h+B���h�9S�Ź�F�.� �ř�{eF����EdL�͙�?*?cu&�/����bآ�������ǩ#t��<|�ߋ'Z/s61��69\�����Q��m���à����y_(�jf��N�]��K�C���j
j�r��&��h1��:w[�6}��ag
��q#�7�v�Z�A|��7�1�Z]��w6"�ʄ�=�b�V�j�E]c^�����`&�͍��
����C � �S
�4$�`���s�bF"����
�b:q=#k����i���w����0.N�:N}�L�Y��E�>F��h\�L~œt����h��k��<0���Y68�=^��1(<I�W׵I��YU�xpc�=�[#���2J���N��gB �)�3n�歆�EJ��j4J�^�lԅVYt��>�-B���9TA�1���?���#n-4���˿�:���C8ro.=��u��5�cN��`��TZ��^'�(98q��d�ZG� ������4�<&�k#��m��X�Ђ�29��K�{y�j+m~y�p:P�/՗��9�ZlEP�=�V����i�����bd_W��'i���ܭ�wy�)�`�!��G������P�d�p��a�3@��x��V
���~����	��^�ؽ:�hҫ��_H��=��$"|���ȍ���/�ThWt��αp
X�~_��]�a!�ͦM������6�x���� .�v綾��~T��m��X��Z������z� �c}}s�w��P�|;��=�5�H���`S��n'���k��@RA��7�;Y�ѯ�w�!��=�Ҙ��(��$eVU��)D��k��n��'��)��qŦ�{%f��X�ђlabj� <M��n������P�'9������� 3y�V�u��B��ȋw��� �v�8�䄍b�滏��#�K[Aض����.�H�{�V��s:2ߟd�C�`�3å9XG��#����3��f��g�7������$3�v��,s���OlO�Ij|;;p/V�ݱ�i����Xg�ڲe���+�NTf���.�BB��&�L0ڷƮ�9o��#�g=<��:\OE��E���I�)�ػ,I�i��ή���Y#�q��!�{T�;Gr�̾�����:��([��Ò~�!�7�{��1��+�)e��FP��ag#�-�ˤ�a��'ٿ�(�R� B��X�Td�d|ePf5҂�Als|`�Y���cО�uݼLP��ē�M���� Z�������t
{�^Py�Gn[��n�ۛV�nU��>�� 4��A�S�>i�����y~�=���gT�|hsl�ȌZ��� k��37��1����*,6�чj&��\uY:$���+OBM�c�SPAt����SކU�m�q,��ފ-�G�&0V���e�
ɳ������b� ��K�>.�VQ�\�"����s	*���_��)�͖b���Ea�:Y���T3��}��m�B��]���x-�X�Z�Q�Q���H3�3�^{��j�m	J-;+m�S5�r��G��˽xb���ǰ1z[g�7�?XC�ɂ��(z�l���	����)Z-{!����L����SZ�v��!�ؚ*&(�3Y�����fT�
3c����@��k���w��#=砡��0���k��(��@
g^�|Ƅ�l<��N-�3F�!SU����fZ� V`7�& �;F�'%������TA��l�Gꦫ�����B�@�f?�܆�=�
�wI7�&�[�ך6�����lP,�4���͔�[H ���9�5�
�{9Ҥ�E+�:�>��;>�N��$+���S����b<�g��ݜ��8㯡w�T!��(�yF��9
��\��T���Y�&�񁲶�i
�rH� ��i�7P�Amfg�;&`��G�Ƙ��à8���~qW�I�x�n���pp�'�< ��D������X@G�C
�z�d=�k?�K�c�*���f��\�_I�:TN&Ϧ�p�����)2M�=�8�e#+BB��{�~d���)�F��#��$�E؞�OQ�K)���:ΉW.�v���PR�>
��m���s幞")j����qr
?9��Mv�N�.��ɢ��|�a=�V��2���U�'4yK�t�t�$������I�U�>��@�@b*|��}KA4UNf4a
\5����⍒~�?�xuX��d�2e]SNȦ�qOC��D{!��l����
����Y:m���M.���L�0�[�7��I��+��t5n㯺��l�>�w0R�ghA�|Lb���n)��9�щ�:�U�H��=i��s�֎0��O�g�8����3��1җ׵R��qB=�*��P.��h�6�S(�a�Ó	����qh Ko��]�����S��'��q���,������(vT���Z�G(�[���7�힄�^���=�.�_������J�7��1\��)�Yb�RHjf[�A`P�!`�\6!��ι=-ǿ-�c�>�b���/��"��� n|p`�{({��`M�@�a�"��n�<��&<�2N�m�J2Y��fnΪ�n12hH��9�ñ�YW[^:E�����Q���d�V�R���D�1w�g����3^��7"�5l��[?���r�y�(�~�#�\�ъ�ln�#�ޣ9`}\C��k����u�:+���_�sN�Ӿ8������V\@LHP��G.spt��i�Mn�U����'�<tQв���G��������a�6���]$�g�oȹ�w��@4~����Do�d�D�u��[�M�J��6��hԹW=`�[��v�����2=��Q3~�^P�� ��3�Q=k��(��.���9�Wj�S�n��.��I^
��!�^�Td� j�#b@���GS@�Y|!�xTPv+ɛb	���_�s���ɬ��]z�`�k�a]�m�^�N�X��0ɠ��N��0�A~�ZJM�ݖ�c�Tᓼ�5$��v����`m:;�!H�MX���(��3�l9�O4c�gy-�.�9��RZ�Y�G*4wc@1������H��)�XMVN0�f"'�U�=��V�,)ŷO�O�����	��T����h�踴�.���qB
r���X�$=���,��cC���Eag���>��PW�?4�$�r.(�ĶZ}���q�75���ƌb%b��!k���lz������n{Y��J�u��f��	 �ȕ��������*�/�wT�!� H��*�u���)��M��a���b�:�]
<�B8��҇���W�d���;W����!�%e~V�1�+��L����� �JYj��$)��6�p�6s�!U�^�|�r��Ζ.���W�h�
|��|H�&�tG�eو�g�0�њ6;h��H�jݥ�D�z �G
�#e�ZZƲ�n�i���8�����15F��Օwo� �>W�X`�� �zu�����P~~�7J��?X���u�Ia�z��r�^3�Z�i����H�S8���H�
�6�ET��W��S�[d}�2)TpfDPK�ʞ��)|ː'N�7Ľ�b�B�y���|@�[�C�7���O�]n�E�b�}� I�F�F�pۺ�����_�,���a�%��6�������W�4�n�P��^���K+u}��f �gX�X�r7��}`K:R&<�M?7K�щ	��#�����4y�� �<��G*$�̩RF%F��]���	�ٰ����ě�)��?ʫXg���R}���U����pr�2�grj�,�u��ؑ��o���\+�LσF�j1BF�`��,�M8��Y�S�Ґ��pE����p҇��\$���nv�]����V�:���	1@�m��޲�Σ8����c3�p�6��9s����m�6D�g�˞3��2c�Ǒ��{���#0j>
�.���4sϓ�8!��e ��	��F����GL�.#��SŤ.�f\�R�?�1)������e9�^	��Y�%'�A�+���u�g��o[�TLhT7~O�c�TΗ��Ň�y;��4��P�2O�r��Kq�h5]��傍�0^#��#�(;�e]e|���%s���ĩk&����g�:�]��p�k���N�Qes>*�6��Z����h��y�$��Yv{��}j�l3tu5�v㑹����0�~	��qKg�����U"M�$÷�_{n=�U���1��c�T�cn�˯vѩsç�"�d𧻓b<���|ب�~Ț���v��T�/�+�-����J�67��������~s ��� 4��������e]�85����0=�S�1�������DQ�`�%ѡ��a|)�%�dh!��!�߁��E�|�%��n�*�M'�*��:�L�UC�T�t�[W}�6��$�o��mlRW͟�ѡY�#�����M4�VP�T��eQ���i�D��O�� $~)��=�	��5� ��6�}Y,����-�t����+����F�IV7~�XJ'��
����sZTlwX��Q<�xo�r	��^��^���C5���p��P�%o�<���.dX��1>28\;�*9ǰ;�7����$�mt�$*��J@����6N_*S�o�M2��#N6� iϓ�/ո��q���l�cOO�L��;S>l'��ni���1��x�K���$䞷�7\�@�W���2�ךt+i��u�*(�<�ĸo� �棅��:
�G�<�CCVVlً�YF$��Y�����,RYEb��s1�Gu@����W������)5Fh0<2��!\~J ��C�������[��16�m������L �M�S���$�:2�ѽ����9����4�q0�e#V�!��XQB^:f��V*��Dp����fJ����k���~���z��� 4��5�|�*�l�iM���r⿟|���/N����x��b}�V�Qi�:�D��R�ù����1&>O���gl�!Q%�K�2�lfK�����-t,����qFɸ��a ��GI��"4��@�{��po ��kHM�ʼ�&fE�E�l���(�|��rL