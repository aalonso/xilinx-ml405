XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������ )�D�&{�N�i$���ܨ�U6�a��^� d+�9�@�$<�C�M��مpSs�#Pvv�Ŷ)� 4C�J[��pabQ]m��G�{]�I��yy��r'U[�w�!T��y�~��P��џ�ivi�a��M��aa�;O��)$����Z����	��'���=�7ٻ�2�)�/��oV]�IyR�zz�Pf|�R(e�x({�X%��cUa\d4f0��zr͙��&���T8F��o��A���4�;��h�{��t���"�
���%"���ޅQ�mw���]��Q�u3�4�
�p��	�<��'�_2Yq��QSsܔ
��f�ߴ��H�J��ҵ�y��=b~J��C��D�t�o�`�������5NR6[�0-����l�X�N�r@77�3�z8dUK+$93�/��}��t��S��b��ZJ��#h5!-�;#8��@?D3���yq�`2�S��������k8� o��Y&
2��~��K�i*DT01�ξ��f�!&���F��pm��Je�-VԳ����b�=QU�W,@j�)�@U������27Vg2��z��I�Igh�N6K8]s���No?��-��k09c����|�iB���4��Xms'*����ٗO��';\�*GW�&�uL�"G~���Ji�sǿڋ-zC�M�XR������9/��R1��ل����v'�w�}%X�g����t�g^&�N[�G7u+v'�|�C,z9d�0;֛�XlxVHYEB    19c6     900΍�����*{�P��M�u	������ �f��N(�4��-VN�~W�_�}��'%Ę�G�A�e���4�6�^k�7?\��gY��+��iˣx�ȭr:�e�aMG#��|��
�9c"����{��h?��\��Ц���L�8�7i2~�\��d�$G���/��Q���Dn6*���Ť�K>�CM����*mU�1��Q8��"���~���6v��ֵ>�Pb�+����������S�m?(��K2�IJT8⵨��|�lՌD�ƃw%XU�Z�.�D���@w��;L��FW�~/W*���/��I^ֿ�nqiV���J�"�i�����6HKT<�(���P�i	�f ����w��h!s��1o_�k�NJ��_E�4�oO����|�?ˀ�θz�4���x(���Y8��u*&g'��x���3���|"qz������ڲp⧤4@�;I��"��b�'8����jL|k��"�9Q�$���;���{�L��CT9|ю %���I�Qrˮ'K��>�m�KZ2gL������ͤ����+��}���W��>�31�淸'����ŝ,���EY���?H.�P�~������]g��?�ٯދx�s����щ�~:-Ǵg�^���g�Om<3��{��G�Q7��sU��O=,PB��Vp�z����(�h ;�@Ձ���yB�F�"4�����経�Pc\�i})��Y�u����h��-ҷ�4����\qڴ�HB��kP�O��G2[y(�����^ԉ���O�͕���n�T�(���y��S�wF-�������A9�k�V~S�1m� A�$���jc2PG��X~Q���|��:��(�K����r��|��������>���nC��6�_�,�����F��ћ`�p�s�p-6����	�_'����6�������Tf�������j���t����ks�O��H�ۥ��Vוt�u.[�]œs��Y�iK�Y�Md���	*�Iq{�40��%�����:)�����ڣC�������*����8��B���Ѧ1(��:���$|�Sy�)�ΠWD��V���˾ `yzJC�߽ �� !�A�nI�\'��d���?�r��._��	zf}n����^���F��]����ց��������v��\���䘼�t�0|
\GZW�uƨb�M���/����#�z(�fxp�,�(kMn,�'�J�i�Ｇ,Qz�	*ʺ`�
�t ���Nfv��a�ɷ9�/ϻ5��\4ˆ�~j.��2.��`�ʅY��k�5l�^@�v����-��v*1fA�J#�{
���z��5���kLKDݪ��wrm��\�Jtjs��C�p^,��2�d��V2Ⱥ�n���5OPSWN���9�t�?�Ꟛ3+˗����xʳ5mL_�!�,/�O�G���b���V�	?�&p�����ޜ��_{�R�s?+����K�Xnw���Kx,���]������>O�����o��Q�{/[1�{]��P���\>ܟ1W @�m^x�cs3me=0B�Mr�H�_t"Q�F�����q4"�Q��i^9���{܂ƞcf�q}�s|�GFE\d[(� ��Ńa�&�!�Lp������m!{��~G�1LjX"Q��x�����&{���Xx���u��f�J�����F�i�lo�HJ�3������d�r�iAc��V���zn�X�	LjM,��[Y�-r�y��~�ϻN�}J�?�8"n	�;��#�#�[�VU+����p=t'2��nUlU6��]�q��.�P��`�)���������]f����V�߾8(�~�lH�y�Ё>�f�s�D���3��&��>��Vc/�5�6�#��U����h��j���My�m�^i�@���%@i���*�Ql���1͕�2#5�S�����V-&3���U�.��+Et��u�A��?8�V�:E���$�v+�ۉ��Y�E���VA��Ui=x���oI�6���+�����p�͝W MӴ�+�FbYAVM���,����:A���:$P����i�lL���6Zb��OUBfT�^4��M�����j�m���^�G�;���װ�?�����;�=��?������p��1lR�+f����(߂ї����f*�b�MP �xF�6Y���|? 6������-�?��̼��(x�C��+�J�"�����X)�l�p�Wth\V��h��vu��n�y�o�c�vg���6v��)�o��/����@