XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F��m�.Eӗb? �������]���?��}����<��������i��t҃�8�=����"}���x�-�!Ɵ7�S���&�?
�4�<"I� i��ߞ�1���}���u�Xr�MW!\>����2��~� +�h�[���In9��V\Ҋ �_D�sQ6͕n�Ę�c��]������|��xX���,�IH���G�*�X~�Eݥu����X�Tی�f�T_4k�����*>"&2７2�������K�E�����[6�\LxQ	����1K,ܕwk�N�����4ii+:��L���������I��R��sI=Ř���U_���W���<Ս��>+Z�>{m	^S��{Wxd��ے�\��j����$#�n��#����Ba�Vן�&	���/xXBQ�O=���+ms�<���l�I��_���h{���4,�bL��có>�+b�+M�_s�K���]��0��w&D�H�+� �0���϶v�S��5����"
u��XXr�!�!;� t����a�������I�V����Ps9�;*�U��
Iò%q���by%�Tk�=
Bi�-,c�>����ػ��ڧ�˸�5vZ�-�K���q%V9�HɊ�:�S�>�P�s	Rs���TKCKH� �n �:W8Y�	����?��}�.�����B>d��LWv+2���y*���v��}>���&,̏��Lq�4W�;���x�S����E�xw����x�km�,{T���XlxVHYEB     f8b     650�Qe�b2��A ğT�"810C���)	T�[�4�U�4����� )tdpU�nF۫+�ȧ@w�דe��;��K[H��5`i�Ar9�~�θ�ܵ�>)��#���!��{o���*��{�b7�PBA�>)����)Ú�0��B+�~+�3��!���5,W�[�^HP�*��G��/�����%���`2�f,}�UR���Tǒ�MⱢ�2"�+�mAP�����:�rs��6�uG��H�3��5�v��9ŕ�Ө����b��F��J��y,$�|d	۾^I��'xp\O6�<tX�Y���c����jꝂ�x6Ӧ�1T/�p��F0w��L5k��E�e9��M��/��yK��K�#��ǩ[�)�����xZ���Ɏ��
�?P4���^UG�esoc��C��n��$$6�A��j,A�����E1�,p� А�_@�7'��!� ����[�)-�挋�zi!~���%aʏ��A���n%CT~�xL�����`�U�pH����l2"G�\3G
U#�)V�����FX�x���'^^P�ށ@n%c�I�1�ɐ�T�#=w�T�
C�5g��l��~eb�i��E��,W5sݧ�j�i�������}�VC��s��M~UZ�B�]���L��}	ه����A�#�wD_׀Qu4-�5�O�U��������jL�	;J�Ev�8��ޜp4 �o�/�a�k[��H�ګ?8��]�����«'\��y�kw�t���t?p���o��̆���Gl�z`ĕg,�f��[�{�s ��ޑU���*j���K}��JV���Vy�����6���ZN�Z��T�k��{-����:�vzFp�X4�ԉ :#�����!�'��,j��6���$��M-$t��n>��u�n�U�r8�/��^[&d�	���Oe"���0h7�����Hdʵ�ۘ(a�Jݒ��05�(d���9']��d�eS��
䧣�er�ꧺB�kZ�w���,��s{�W_J��
��v����2�	��̮�H�5�?��`~�{��M���xY��>ZЊ�`�����}6��שV��Dh�h�l��;��b�橥��BO>�R���ݸ�����~][h'`߂�W��,����-���[ܠ�/��)JY��Bm9{�t��<��:�∆�"��&�E#3;�|S��o�$ ��ꝷ/A�{G&�0[.'O�v��)��X�	X޸�������b|���{wИ�

B��Ps�2@��Z��7yYY�}Щ��U3����>|~,2Es�):��[3�`ؔ�7a�N�Ln�_j�eF���q�ΑT�:6�8"�qtmp���F�)���w��-M�a�hNc	���M��~-��R]��Ԇ�R�-C��lVX��'��3�C<����[��]ڻ�{B�l�k��w�Tu�}�}R�_�2�9�����5~���I���1FxD�[h�K��Gg�P�=ϟ%�}t�1[����`Èd"ډӂjh9h�}KL��K&���$m/�?���ėrF�S�?4T'�wC�:8��u�w� �)�9���u�����C��Z�m�E{s�.#���2�8�m�&�