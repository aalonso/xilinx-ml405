XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1��8���t�rgOh��P̼џC.�Y��*z{z��S�ȹ�5�K�b�-⌣Ɣ�<�B��(1.f]������������NJ�~Z�ɮ�]7���ؚ����Mu�p���L66��;Y@�Y�Z�N�Bxȝ���� "k�B��MY���˿Tڀr31;��>gC�19��	�eP%�/��>���)������6��:������ɛ��GL���.���A���D�qe��	���V�);���C�����j��h]���/*#k�+	Jm��GC�B2�{��Q����˞�&�������"��U{��p�Q=�[�\��L�J�Ϩ8l��+�h�����J�Z,n?�FB/W���j�g�����$+�.�K�
��9(��
��j��`f���/��N�$���%�e�dn���$�����h��ٻ���9gE�
��o�`�ۇ̉u���.��HW�`��������Ƒ�	�8cM=���s��{�����Ӽ����pK�θbK�|�8��ҵ��X���&�/iq�d;�\h�`T�sa]X�^�����ף5������������ҺA��P�����ax�:A���G|]	B&�ao�����n]%���ssW}����L��9�^Ͷu��tjy+F��0����5�$ye }wF����q��3ߕ��. ��ƕ
�y��q<c�ѯz�'�:��{(�JL>n$���v=����f��5�u`���}�f�f�����Y>����@��*fXlxVHYEB    1661     760T\Wpm5Ҟ@��������\�?��7���:���Y_�_���E�(�ʷ�����
�_�����"��3���\��&o��S�m�dr&'���ֆ�X��,�Z�` W:���Mv��r+����CǷ'=�ݶ�˂��F�P�a!��W����l����za|���˕��mh�W��d����F
��(���;��ߒ�x��8�5M诧~�_��X'o&K;i��㉑��ࡐJI��9�@޺����3�gV���Q� (��>MY�}�3:�7�,f{�\-��p�7�
9G��g��H���l�	��iiJ�~�I���1�E�sË[3�="/-�XI-��d����>�����E����MT���#��ۧh���+z C�	g��i�/�[4t7Z����ٰ��?��J\;���1��+ȑ7W��z����y2�T����r��8��?�^��C�K`�9�Xw�O7�9��������0�F.����]���s�Po�ڄL>^�����k���$# � ���"�=G��'>�+.7�m����,Z���T�vk��h�i�Xg�C]d�cd֎Z8�cH ��U��Ry�c�$�����0�/�ؚ�!�;$cHFƋ�_Ja"�T����YG'Y	[w$,Խp�j�4��QΏ��uY�S?��\U���ox�s�:�8�O�="-u�v�&�a~V���pp@vO^ƥ�W�\�zt�Ѝ�x��k�f%Ɨ��g�@Zy"�8>����Tw��A~��>��)j�>�AU�N�|ۂ��j�7^Y��M�|~�|���K��I6˭��^��<Ho0�=F�%�Y�D�C�JQ>�F.�t����Lߔ�TI�d!����gy�Om�Q�62����(��`1Qv�A%�/tʏ
ii72���������w�U�r%����:��0`���{:���M�9�thY�v3�-�I�� R^P1�7L����lLo�R��P��T��}�$
���'���5)��ʦg�C��7�H�]�<m��j���5��Л��dT��D��r@ɜے�~T���Z�XH��LΈ�%���e����@��bG),).��C��>�=��4A/c;�W'l���٧�>n0�P�X��)�Hlq�l���G�K*����w��/R�t�Z+~�Kw� �x���������J�Ƭ��iv�l^�(�El��Z4e�P`��� ��+�6~DMYԍ6�c��=/#��M��<T�睒�^?�St�[?�v�R�<ш�<�g���(y��3�D�9j��q�y�UTN��$�9�$��}�b�{������N�����	#*F,Aiz|����g���e�D�U�L#�IU���/I��ӏ�m��M՚ٷ�Џ�`�3UV��G!`C��}�����
Ve��Vv@��{�+���^�*[Q�)�`�*"^��$a2�Zn�U���ӄ�;_�8'�jX��V�{��8|>�L�$�|
�eE3�ur��r�v+��x����ݭ�Ÿ<	��m���|R!$傒`��|kGǶ�8�C�t��5����U���Ucլ}طg��:I-IMؠ!]�d"[ȸ֍���
TS8 ���S;/b!}\R�-	���ױ0��ܱ7:�^�sT��Ú�j��[���������E)�jDva�$y���y�sSS�A[�v:ޭ·5G�W̿|���Ӗ)��[��!�<���i��A�mT*T?yF�PQ��˪wJ)O���hF�+�D�v�!���� `�����h�rS߁[syή~�$��ڄ��`߯;�^�To��!X���+����g����F5��E��*J�����#��L��&��J�QX	�%+�Ҽ�f~g