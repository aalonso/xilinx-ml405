XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(Nʹrz�a,����:���l&��17��i���leH"d��W��sd�_#9����?K�P�,m�C�f�\�ʼ N�G���D���We�5��qR]"�`0�/AIM�+���E%:�s�:�'/�<�x�-�T^L�G��-j)4���7�[�:�-�2!,1���a���Pn2wFp�2�����Ŧ!��8������� /e��.[_-�kX�9��l�V[ŋz�B���6��S+-�*7W=kzC�{7�EA:r�^�w*>Y�(Y?��w<�]5�z�q�cM��Q�r]���?��V�Q�����`*���a:Fd�sg��}�C_��ө��*�).����
6Ӎ:Ӫ��ȷ�>X$|��G�`-��7e��jH��O߸���(ҕ(!�E S}n�P+���"�T��æd�ffI.J$+}L��AGlB4�-�|qk7ِ�,w����\{ �<^�{�Y��w�C���^p�B�{0�M9ֶ6������]��0e�����x����j-�Ǆ����%�QW3�[+Ƣޫ<�QGp�9����І�Q���]6��ǅ��}>H<������:���XQ�y�P��t�"S�[y��lep5\h��}?F�֞b_�3�d�q�Mmn� ��@z����W=L_xJ�Vȗ��_���%�Ie�o1�R�1�>�cdv{�����\Ⱥ2���4�-XR�O=n^]8�`(�VU&��n�P�RQ?�J�2���'�)�����z�����32�n�kQ��.�=�9#n+>�W�SVXlxVHYEB    1111     710v��g�]�w�)WB���D��N㽵����ɛ�,�fF�ND�9���-���!�beXC*8_D���0s����Q�Uֶ��c��<(M�)�o�\��B�e�R�9��?O(��hx��훩����\(0���Iё��|F���$άW3�Yy�#=odhK�wfW�-[�BC{�i�Ukc�"-D� ��T�C�RT��ˆ��G@uY�ݜ�㡽'X�.�s�~�I�� �w��hh�uG��$��V;����{u1������n��햓U�E�G�5��Ű��F�#���=~�Ҝ\:��/�i�Zz��FA���.Fů�Qf�*0p�I��QB�D�����b���^���^���q�K����i44U��7C|��~?��7*eg̞|
��\r+�p\=?+e2���}&���%x,�[�|��E��I�� T��?9Q�����9�ВzW��8����)����
Q���9�o6�]4`�sÎ8�%.�k�j%n�*0����A�*�]�s
��Y�5�kt�������r�}@%0��0���V���mR��z� ��O!�n�"�T��,���w��?B��7x���,FK$2b��vZ�^���]Ȝ{(y�&h��u՟AݢW��<�N>|��dH�~%,�9����Ʀ�H;����[B�ƐK�=Y��+r1<���bo$�}�/@�`ud��m�ぜ��ăcj�{s��!.+����$��ɛz��j����M��D���)�d0s�s:��p���������N�Qrڠz
@���!���~t������N)n�Y����T�_h-Q�N�y�h��.�p�W�U��!U���PϗYc��&��y�6�vrLT�y�S��^n��5�h���-w��=0��t0��I�d�-=�F@\Y�<˹�vi�uj������pꭃ��%t�pf��� c޵�����-���h�R
0�i4p ����4I�X�/_@������iټv��$S��Ԓ�"��p����)��;�ҎІ���Y2��Ә^M��U�ߍ���l��kKbu�p��{/�O��	�Z�u��j�Z��Y��L'�N�+}o��[�`?��O]�����0.�!��N�K�ꕔ-�
J�8�{j�� ������JЭ6�!�V�O�̬*��2�0��$u�N��#k��S�%�n�}��g+���-Ly��=�~���M!8�a륧�M��r��
�����8=��`�t�1|�1�i���9|�,�����u���Ȋ;Qa[���3�	*�طf�~���1���� �w�9�e�7;�n�	R�1[V��)d ����`�>ґ��"o-�Q��p�+魐�Y�P>s�=���v�y���3i�%j��T��g_���c w�G������'�Ԉ6T[D׀��4>�P���YO���)k 5���Ү#�g���p�Il�:߯���e��x��<���͟��ǷvM��9wj����^ކ�P������y��v��wB��
W�;*-��T����6���R�O�oć1��'0b�i�fM*��Y �P���B "���P���SEи�^y�f��'�R5���:����3��WYċ7���OI\`�����ɔ�H*�S:�fg��'�Y��>hsD� ֯�hB;C�~�9��#��r>3 �+b�66�Qӹқ����G�Ԯ�yax�'����1��o��vH�<�YC��z3p�9�@惱�Z�F��� ����d!�$��Y{�Vf\���t-�΂ȼ�0