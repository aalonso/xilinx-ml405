XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���.�X��!�*p9���
�j�w����Z�h5ks9��V0ؠ`�F�ܪc;zk��_�!�}�5]@m�!�0�a9�H�*��ds,zT�?d�H� u�o�+I&�è��؅�����k�p���,�J�6����(� � 	�8(�[)l^����X�������~��j�Pqo����/��E�%��{�dw������,�!�Ɩ��L�ո�x�Ӥ�Տ,K��!p�g2ݫv��\�r[�\p	y��j_���j�4a��v+b�ۋ�Q�E0�a��%��5�t��7H3o,��i����jM�f/|��c7�$��<��~�I`yڕ���ޜQu�|��� Pq5�x�wֽzw0��$'Yߛ�u~	)U�0��0��Z�_�+�Oi��W;]fN5-;�Vl2�'|�"��}�i����v�8�]]_��1����(O�r�+�%��j�.�.��iV��c!Y���+cb� ��cW&�A�,��T�,�	�>g�?�1>�;����q�B�����i-5q�Z�� ������1�q@6�)��o�	��V�+!��u�V�j�,E9Y#q�5~O_O�4�g��kRc���¢~��������������gVK��hۧSe l̹E-���zi����\��6�p! �v��K����ՁM�8_/�>/\�ռ �}���m\R<}ó^��	ET�íl��{�U��1}���ٝ�2}r�v�ע�,��܁��~-����L�V,�<�n��������uP�6pxXlxVHYEB    1854     8a0�A���&v�v�0ݙr�s��UD��)���
.9��~ M����,0�R��B��3�(���>���F�W9�L�cX��] )ٺ�H��g��}j]�s���D�Z�?�R{)Onx�r�6�}���9r�p�PKN,�c�$���z�������,�:eS�.dtw�5�F]�D��9q�P��1ٜ��mIe�?�Y�RV��R�W��i�d a��-zS���������Մ{��X�!��Qh�� ����Ei+�7�cU
]���H�rn�	����Ba���c����dGdn��-6����v�n瀘(��faV<�5.`�8q����=���+K3��;�3w�njT``�YH_���*�w�m�nR��6�;}'TҨ�!�xAْ��{T�ƾQ=������ܗd8m�9	���\���d�8�cO�!掛��eI���x_Ox;I�=Z(L���$`wJ�/�j�Pb�H����P*<N��%Ę�5�:M���+Bb1C��������RW瘷�}W��G�F�6���y+���E�þa����6��C���\�s�#A|�O�1,���3��]���z������V8�u��T@�l��d�Za�3".E�g�d�$sIχŝ��E��̎tzs@�l��U�'�KG;����b����4���^zu�4������3���lmo3&�`�2e�a4Z����ɆCO��H)�F�/MH��`�vuv~�C��*�z��(^�@����#j�u�j�'JJ3��x�eK�����Fa���d����F;& �$݉f@�X^�> -�����^���U)��ŏ�ۣ5u1�	�{����uLQ���ix�>����pHe00
8�5��G23��T�>�bZ�;[e���E��pl�kp� �LH#���,��ՋD�s���u�
�z��V�cއ�&�hĨ$�R����-л�7YǺ6�k���xvc��x��Q��6z�ýF�5����a�͘�>!
Q�4I/��&ZT̃���̓���}r�V�V��pBDy��&m�!�5����g+mBl�?��H���E�7BV>voa��=����y���'����ᑷt��sQ��e�Ȅ-絚-�p-�r�C{�=يʠU_��~�W"ISZ��I�U�!���{��L����3N}%4ì��BE���=ݙ-�-i�����I���QL�q��&C��d� ���e�g��#��!��u�g�`���9���e�f��-L�֌��c�NV��E�G*Ks��v��K&x� n�C����`�5}��h�|�֫�;�x~��*��[����]�#�6��,�^�1dnnb|�\X�i4�5H�;���y(��y|u�Ma�Y�^LBj��Nߗ��U��� T�_TH_h�������������/u<{�Ě��I7�`��`Rڌ�M��QB*[�>kޕ��3��S�'B��gI��l̪�;rGx���H�	i�䗲t�&���^>�� '�Z3��,�1�r��{8����a��yO��y�S���ł�VK��=�9�8;
�⤷���N���F��p�:��<Ma%�RȨz��Ѐ�}����:���!en"LR��c1o�q�?^��$8���F��/8wp�Mi��Ӫ�Xc���tEowj`�]�}�S��$V��\�%������4d���ey��;��JQP'kㆬ�R�P���!�?E����u�_;d����?��\Ƒ�KF7`���"���!v:�����
�_L��%���F�~6�a��(��+��-uP�4"���R0�)b(X`W����#��
;Lɻ�U�������\ձa I�`��-�f�5-'���W�CY���b��:�&�o��*%<��Kp/��0o�@(,4Lg�]8��B)#	Q0UF˗��k�ܷ{ҟYč�u$�I&<�)�Cz��B�W�X�+#����˘�&��2E���TJ�G5}��X��Zi2k�e(�Vׯɗ�Y~ͽ�t�\��k��.3�Kh
���~ƙ��Gf�E��E�����e��!ʚ��+2�~M`�3V�t�� �GT��Ş���31��m�Q�P���n��%������Zm-�,?�<��|��T�X�+�5�B���'=o^ �*�n�t�q1�;��~c_S�5؍�΢g�w�5�@ ��b<2v�G�G�0�o�.���M�U�