XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��XFƕ�q��3��r/eg��<B��x^�.;������U����)�7x9�&-�oNH�[�Y�|&4���H��~ �WJ�RsH+C)NQ[��dd߼G���x"rB<-����S����%�wR`Ռ��W`1�,��c嫰Fﱶp�Q��/r�'��g_:�	�&�� �I� �M_�5�����vLk�W��h�Bx����aGR%f�mJ�/�8��bh�O�=C�펄��"�,v����d��V�P:�h�ޯ���)�_�}���Bg���hO�n���<�.(o0ڈa�d��%��(�Hޅ���{Rz�0�]��j�E������4#���`F���Lbms�W庡8�7����$
��T�ߙ�,�Q9s�,���RÛ�Q��Z&��fO�K������*S;.��T�n�b�s�k��.cwy�;z�#������ b�{������]�Q��������R�!�%�x�dR+ ��ҡ�8'N8�����\֗/׍Øh��R���=.��g���v�����wr�ʱ;o�����2�F`z��vr(�i���a8�7;���"�S8	U���w�6+iz�lh��<r���g�Hu����x��3�"�a���|6��V�*^��Fm��������C��t�-y9N^��'!�.&CԱ�[B�/g�I;
*��t�A�O��	ԡT�Y< ���J��˃ԫ!;�-|ۮ9>Ã!�h�֫g ����o��L��y4R��e<� c�%s1��V�����l�0��8�2\�����%���v���AXlxVHYEB    1d01     a20F-�z%.M���cB���]�o#�1��g ,��8O1MQ*x"ȋ|m�wxFn�>�`���f)]x]�s<I��íݟ$�HmHp�i�e`:�tCW�lc�Po��I�(���u:���q���,�+DHT!@���6oy,�'��,wj=¾Z�D�a�>�FX$ƗDʡB���u4�1�g��l=w.<� ([�]F����T*^(�C/9w�]jNsx��Ӭi��.dm��iji�u67\� v��2�W1MnP3�j�N:>l�`3���r��?��Ux[zX���&��d�?��,&�#έ1�5�D0�S?��� ���a\W:/OE��ٹn���+��%K����v�1�!!d���i1j:id�e��/afD���M��3&�mh�Ih�d�슞����t�^=e�e�����K0^ɍKV��O4�l��j�X��n��Y]��W�r��,B�rZ
mq@�4�N�Į���i��A��{��絊��kg��܆{>M=fp����l�gxU���%?\�ן�m2	)��Ná�l���\�}z���cۣ��\>AP�AW��O� v@�#�Hq���mp��OQ_,�<.��ܩ��#�1[JW�2���AzUt��A�h�p�,*L�����.�`���u���Y�b̝�GÃ�it�܈F���E��2�jY��	x���eu�-�K'����f���@Y��cY��k�͡�<`��Q[��ެ6��̌�+b"�a�	W�3~֣8���::�nk���O�r��f_a��j�>SL��<��.K���,�����j�U|�6�!ao�vQD��~9�+#�I��7�4�MM�)@�PqBV��I��xVQIgks���O�s�I(A�7���0�X�w�! �Iy���7-e������ӳ7#�k��܇��d���ޢ���9��O�;3�#ڥX>$��p��]�)��J���O�������`]�V��s�<�}��!j^Y�p(|��d �����k���������cg��x�����uqvVhL�F���1�sN_�UË+Bm�3��f#�}���\q�WI1���VM��X�u��؅0�d�)ބ��^2�t��NO�LP����}l�!�b����k��k�^���T}���)��S�5�0Ԭ=�>��C�3P����+����Ҳ�����}�%�7��e8�،�j���p�N9~[Tj�AmY�0;�A���0,��иt����6K�Z�z�`x��S�1�gN� ��_	���0�^9^7��u�q���L�:u�n��=��8�]͠��	���s�(7�G$%!w��CF�KA�� ����cj�-�t9��Bu�..4����J$OLCJ��!]����{�}���]���:>�|�hJ��"�J�s	������2/�ψ���R�����tY(#u���S^�J��;���>!�g��24��y����KoX|Z�WX8�3���F��`�Q�F�d����g+.�h�Ms�ї\E���}�F��R~���sm�ݸ�	H>賈�Z)�޴� PEd�~v{k�x��AۿV�&iow��=�~Y�@�l��/AZ�M&i��g��M�<mRZC?\�k�$յ&�x��8�TT���`�+��0�Q���,�m���峝��}�dsd��	g��8��2�L.�"��]!7���z�R�
(��e)�r��
=���3�샚(�FrP�r��V��C��7z,I"���س�^1L��C�N�V���e���P�\Xm���≗��`<0�$T.cU���Q�:Y��$���y�1�cU��Y��lk4�o�\W��l�ݣ;�el�,Xl����T��-��u����'h�߽y^Y�
UX�n��>;
��)��aM|w0���_���0^�3�1+�ΐ����':>/����:}����<4�Dt�Ţ���rCt�5�!�&-����b�T�Qq ��{D�f�7̮�⾘��H�zQ����G��j@T �ޟ��|�j��;T������%���s��9�x�M�e��ϒT/��?ז�}u��޵J��lO�����
�\������Jd�c:W��І/ktIL2��%N��b�`�OQj�u���	�X�3�(�uDa��x6ő�cR�{�*H�	I
��ɲ"�IL�0��h�MR�b��-@�7� &��gv�w�ȒBʒ��[\e��R5���Z��9LM�s�R��:���q�y� #,�ukd��s�S��다��v���I��!�9��'J�"�*d�;R�D��?�n��;��p�g+����c��ܴ
� <i<���~�Y<�ld��l��y'�\�9�\�"3�j�<���bxR�'����k�W�1L��S�f�?٨a�e5�"=�gIOk�l6�ˈ�#���Q���TK�A���۬��G5-)�at���WAY�� ����������c�2Igo�("�j�^�,�ft��/o lgG�����1�PW-38��L�q�C6� ���P