XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&r�+�6��2����;�[9�:)�R��Q,k=�b�7��9��xu��
q l�Ǽ�^���� �aN*�8���b!k�u��DOF&!`�AH��������+��闞f��ۤs����gBJ$�L���i�iYG�Բ��!��:�p��rf[X�2s��%����fǠP���Z�s��!VP�*Z*�rK���ʳ�ШN^z�[�u�<��W�ŭD6�md��D�|i_4I�mm�����.��_�P���X��tC#��"?QEBj��=����$�P��m�(B�K�t����݌�^/�얯��u�`_��tk�&z��<j?yu��۝ZĥV�:}d p4�i�g*㝃�L�`�����K��x�y��c@�È��%����8��6"�Y��ەj��M�P��'�ԘT�#.�L�gm�i���z�A�R�t<:L�mef�"M��"~��kO�˜k�8���Q(�
ңn�OSJ]�g�>k/w'y �r�Ņ�o�fǼ��3:�%줵��V|J�G���$\EW�m���:��#��ڡy
�QU촤H�4�m4CPPH�(*|m���N�u
�MIxM0�}�Ӗ�9Ie|�+R׊�px��PrGc�V�!ǅ!�t��$�t��o�O��jׇ� �|(_�o['���z]�"�	wt@��DC���`������5��&�.���#�Qg��"���2,�%���jI�pG�Ё�|��a���v>jNnĂwY妯����u8pr%ǝ[����XlxVHYEB    2fbd     d20�,�r�݋�D�	9��+��N�-o�k�I��;"�V	Ϛ��Jv8�s�N˖�"���׏�}��!S�}���J�pe����E�LF��#��g煃�v&y����rq~o��̓N4nY<H!��4����<~Y=�a$�M
1�c��^sL1i��v�bD�Ygᩐۄ�^�`O�W�7-ZDf�%�-$�Ǯ�Ԍ�b��=Jg�Ay˳?%�7Il�� x�Zt
	?Y0� p���i1_��U����7�O!wT����\%~�E�_#��o��٨��L]�Y��Q�ߒ5���wܝjG�G��v�����"�<P��z�j5��4G����r�ȏU+/%
�O�|�c�!2��V�sge����	#�<�u�y��\Mb�=��Vm����8��z@��;�ή���i��0Y�n�.	�ǥQ�L`۝+7���}fg�e������i2W�w��Cl�05JyK��c���G�a�w#�D�_�
H]�}Y��B�7E����h��%�0�����E��?��7P������g�F���_"�0�G���g�ʜv�tkI���JG��V��d5?Χ�4��f�Ύ�3�
��
Գ��a�-Ld8K1f�ο��&�������=^b,~�v�U�c�ɿ��#�A�Ϝ���/����7k�+&��m��Ϗ��nl��6��ruԱG~���ڥ]����w�o<.��
?���snY7Jc�\��������
��sTΒ��sӱ�j7��L p��v�Q'H��e񝶌�8QCE�B2;ء�C��TǗ����3�JV�be�"�n���	�)w�'-��Wt�x]�m��Oy�����fRۋR|59EpYƤZꙝJ�5f�Gc���kK� ���=�|},�u?�ª.��qOY%��+��'~~��%9��ލP����(��,c�@Dp��{�=m�n�3vs� )d����
aɗ
�)�-��Z�Wv��eЛ+#�j��S� ��B��3�\����&��Bč]y�����k�������BO��g|?w�Y�	@_)-�F�$��-�C�"8/��a�0'<��:���#�(��V�P3���ψ���+����dƇ|q�W�0FW��2���Ee��3r-���ny���O����[��
����Pw��"�Q�1=J	����
6�6�*m���W�\�_\fGUΩB������|t˥m���TMm�"3=�y��QJ�})�w�y����ˀ$��a6�i'�ک&Kb�OH�~�a��=%g1��|g�����	��N�!o *��^Pv�}�������E��(�rA=gU�J�����kqи���]ӌe��9׏�/7(���=9��7X����,>V25�h,�:m�@��qF>{,Z{J�eqG��s��y%��s�����ā�n���6s`oXC�x���<�a<��^GJw��������ǃ�8^Qc �_\�u�g���*�C�\�3��׌�F�� �|͝^���K������ya��m�"
~�9d)Gg�^�f��3��g��%���X���hӇ`�`��՝}^�H�%��ٕ����ys�ޚ���|�Q'���0RLU�����H)+p�����k�F��Χ�(�Y�R�V�4m&�wL�����z�lNV�.Ͼ<�}U	�1��RVx���N�2m ;$c�֟:�մTP�ꮢ�9��g��KƢ�K��P�L���:��|���I�[�������Iupd[4���s���fJQs�����B�)-��g�%��������C08��u߽J;n6=�'8DoLn�5^祅K����@,�ϓZ��&1τmM���7�Iѡ��#e�y���A�gS�@CH=��V��`���4�~���N@S�<�JeY�A&,z<�<��6�k���� �"�"�w�_�&;((� �)�B��7T�dى�V��%tj�Pv�*l0
��U<�IYg�K���s�n?k
����a�Pn7(x)�]�Ux�i\�Q�v�U�#^#)�HYB|.eu����X�s�=�_6]y; ���S�"�g�t~�!��N(JO<g|R{�n�^�ނ�3�hU2�T��Z���.���_��՛�iSt~�nT_3Z^�˰<�҉�Ev�=17���"VAI��<���C�_����T�޸<�.�N8����:�#�'����p}�R�3Y~�x����!&��_�/��-l!:�z0ɺ؛-)��̙�î6�Oe����|���&�!�ͺ&*�w���,�\ |'�ԓT�!����磍��z��/�|��ⅴ�jz�\��K̤}��������9�K��rD�`��n��n�:��KW"��������(`�z�,�w7�f�V(�MZ�m�<��-��?5X��xpYkŞ���)���?U�um��[�T�J��i4p(?�E�"T%���<�"�U	��9����\^G�����5p�WL�̣�ƃ2J����,�����c�)w6��i����ooܙK��k1Em�{DОB����y���qA�����G#̋�0 �k���7
�B�G��q�Sy_9Q���n�߄���i�Ɩ�9o��R�U-��Q;}���պ��v�jg*��v�$܇�ױn��pgGC|���h�L�M}/��hɅ$T��h�"��A�D�G�3!nz]5�A���/df��wQ����_s��ۅ�!nx��q��'^GF��ܖ��<Q���^t`��n.��-n>Qe
"�9��h�.W�i��~+�����,�o�A(��|��th��0��]��x�jQ�RQ�58��&I��]�ao1�@Ɏ�cj�QH�����}��S��(����0�
�c+�~�o-e��g���+)��?U\�{���Qe��f�(�Ҍ�W��M=�����x���$Q�G�������ة#�?X	R��J�y�ElXy(S���I��_�DthW�D]�c:�aN%�`�d쪲�[A��x˵�ȩ��Tax���k;�[�2>�[�����R��k�aX�15�J�����p6����Vg��
|���nY�@"զ|��c�$d�[�"�mI��}�y8��{�9�r��eoWP��c����;Q�C�.9=-)�/є�S;�$�)�L�8�%��?I/�WI�2B���i�����#r��J��z˃KP4���3�r+lbu���p\	��G�`TҪ��wN+��xҚݲ�e�>V���(?կҭ$$K������ٍ��=��pD�����oCM�\ �1�Mrh��x%�3:z�Q�z����7���.v|c���p�|���&O��mb�z	�^��!5mERH��MA:xߊ��b�#�