XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����F��|�P��3��Y��4�dG��]F�z��#"t �u�n��s��:;K�V�t6�Yo$/C*�b8&	8$���ib��������QZwK2BS]�Y�iby��1KM��,�Tִ���7B�P^�[h����!�Ԁ7N�.)���O�0�٩e��o�y��.tW�,%`�H�i��°���>n,M�����G�����H�ܽ�Z���i�R#�=x���KBK�/7r)���3���P�%����������j������5���)�d��w�?;J
7\�C��*J]OR%2\z�8Iө�� ���3�_���B�m�ebL��̀6�=0��۝ף�B�̡�ML��q �Փ�]|IU�q���**7�B�\��{��e#m�lZ�:i������Q��R~��X)�vzͯp��	E�� ���0��q7����n4I�폊�s}�'��܆�}Ny�۷���)�G�8����x`5�	I����=��Lܒ�:V��N����f�`Cǂ��P�Zdb:��S�"�Z�

�v��{��Y: �x��Α3o�Ի*R5�]�}��叓[������`��+���$��z��a�%� ��Yt�Dy��Rc'+������_!;���K�l�+T�P��~��V��⣺�h�{��p��A2����$4u�jA�㏖�`kO@4#1��%���3v�-CU)a�N�w�!��=������*�kfL!X��40���XlxVHYEB    1a2b     8f0���B���B������gbCw��Vi��z���p��s�1���~,�6�����8
�|�#�5Y��s�4n���Ф2a�/@��� #�$��y<���r��D�s({�^��s8,4����^����~]r�+��74���,{A֒!�*�6��`|��o�Y��p�����+�Z�˾2�s^�E�r����K�e��86�/�VB��8�����.����c� X;��g̀�!G�^&_\��,:�lɂ}�z�i�q��"�,"��Id��t�.�\��SP�zi[9lA{J{_SQ\6���η�dO[G�Jc�Fx������Z�W��x��W�۷DX�>���2
�y[_��h���t�͖���+|�ML��A�J��`(�v�So0��B���T���]
��-�U�!�� �3(ƪN�����9$�1<,�Z��F#�GԹh�.�d�%'�&˽��!�:�H�ʹ�Wn�� ��7��77^��F�����F������v�۬�rA��o�dp�Ջ`u��nz���&1����J��*�W�h~-�
B��hV�ͳ��4�0�� ��\��H����;��`j�������7��Iڨ�L�ۘr�rDq7��o���U���~U�5�B��U���L+��pՓ�w�u>�j||A>U�ɾX���7a�im�jY8���#�V�_�0���\Ж_�ˉ"�zՋ &u�-��mP����\���Z~��t�"K'�.���w���f�(}�ʔ{ۃ�C0tm$��h������q���v�'m2OP��k�>�5�Α#}�<����Q����E�t3☆�p|�eO��3��l�����J� ���R\w!��8�	�_��?	���^i_v��t�
M,��*wmU���-�H �	5(�d���UR��g���3B��oD2G��E3z�[^J�Z���ld��}M���L�qN|�	�H^,�P�-.��t�ӻ��$x"䛪 $��$H����2�y9L�/�M��w���uӽ��\f
E<=y5Ŕw����S�I�-	�� i*�p7hW�%�?.Wv���/��!'W� g�_���#y�:.�A�0�`%_�}�Mĸ����A���Ό�ؖG�-ݗ<���u��+�@��M��y^䡩\c��
�_��A��~�4��*��b=}��4rV�(�,J60?�[�n��C��<䰺)Tí�̽jH�c�YV�d�=(zu�ke��C��,�ȗ��,>��Y/H� ;�@I�SJ��M�-L��$�bݾ[���� !$s4���V-��D��U����NA��e<��<gRŞ-z#Sў\�,���]H�%g	R�C�ݖ���mtY�%Bų�GԨݛ�����g,Bp�j?�<z�y��l_��r6�Ut�2y���s9^�(8�'�}���K)(��e��]�twQ��B��-��3 zcO�t�g��@,���b�����b�D�f�|�S�D� �&qt܃�����&�Cp��ޥ������Gָ@BwE��wۣ���vuY	O������#�gvUY��T��/�J�I�N� %���D�k31�5%��RF�W��c�d��JF�cG�Ȕ�Ș��;~�6C�j�(%nr��̒����nՊ3���oȃ�qf�@U#�SZ3���E bt��w�kF��/�� �����-z�Y՛*N�l�V��Z��x�Wǽ/�V	5��0b�E�E<�6I���o�4~��q���BeE�e4|�8��1�[w���v�*�(.�kYmf�p����u�@&<�#�7H��\�`���O�KS��H�>����.���?��vg�F���Qy���=2�%���+Ew�#"����a���
Tݶ��v�ue�)����2��@&UZ�_~΀&���oT�[!XO(|��H�;Jh$j'��[��^`$�,y������
`O�(�V�=�&@��v��A"���oQ�*հ\�F�JHʫQ�^�V(���z�q8'����^���`����˅����Kz�]�y�{�����̟YJ���G�Ȍ\���W�̚^i��69�A�^�*�i}�|>��m;�a��a��+㦫�)Lu2o�0ܨ��p-�%�?=6�=`:���Y>�����CLv�����@��o]?=V'j�/��N��B�x��ޝ|la_�9ͼK��D�8M�}�������2�������/Qεm8�i�;c~��cD_�!2s(��q�c�,