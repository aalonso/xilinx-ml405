XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���V	r�7^����6����˱�=v���lr]�	��4�u)䋩�'�w���bW�ߞׄxZ����w��æ%A�1�,�.�i��T'm������N��i:��2�k�q���g��v�~Icle��ki�5���|ҿ�0�Y����(��(�T����ϝj�p��1;J:��ދO��t�'q���| �Ɏ��֋ R�����9�J���;C{�27!(�(�݆����@P�n�QI"��P�mFA\J��]�63��g�����Mh�q%��{�9��^�*�-Rl���c�)��*ӏS�����A�Gm� M�vD�H�l숌^=��P�60!h��c/%c�|t�n��]K�v���s5�{\�%�c�F5,�4Z2�� Ʃ�$h�0V��;u��7�4�9�Q��ʺ��#���~Kf�+�J}��"eگv�B�*W�0����K�2Z!>�X����I�Ĩ�c/+���#zL���"f-�jmT�o?7Cf���A�F<�3��`32qU`�ԸZ�t�^�g]�ijN��#g��FOM�����¤x�V��
B/��VM��v�ʼ�������'1WW����7߆���Ҽ��}��'6�����bM�A���~�;��)<�?=:�kע*
*���|$W�܋G6�g?����O���֟Zlc���O�2�����eT�U#�fA����Q����U�,�\�Q�q�_�2#��*u�[��2eD����9S�e�o�!�q<#�L_ŕ}շ��J/}XlxVHYEB    5f5a    14906rX&����kl���,���k���g���fŗ}����@�h�!�-�Ȧ�x9���k�/��k�m����bl;��ł�j`�,\����f񂌗�7����x�`�H��[4 �L�x�җN��d�E�}�ݲ�4��'U1�m�N�����|YRoh���4�YvE��9�7�n���~.;�b�Yq0��D��}	����Z���Ƽ/Y��P���s�����[��[�1*l����U���b�ykM��_�r᫏`�I�9��Q\T�`]DiJ>y�0�:�<p���j�$)����v.��U�{1?M�&�gq��#�b��7x���I�ax(�82�������\�L�M]q+lB��L�#7v���-��������X0 A���a��g�Ll͵�t���X�c�H9d#:k[����F�F�oլ�Qd�af2`�/�HV=�0�h�j��4Q�ʕ~�FK�众�WW�|���⻁'1E{s,o��������DD�Ej1:�����J���@�����+�
N
�j�� �����Z&(�*�\Ej^����9I���{�*ϺX�~E+�>T)��C�3sVEx�(�f7.RO�y1�GcZ��$���6�s�"DN?O�N��D,�tZ�-�l�f�i�l�hlLN�ӊ�i��-��K@��ң`ظ�d��g@kZ�Aiy�	��4�._���l�S�#�j4�xf���j d�40�۠�p&v����w53����|F`t��l�q��(V����e�
<G�B��9��H�]���+���E�_�[�Rn���nB�0H*����$�DDC��?��_?���:Ih��R�(�1�4��d�i�&��(h�6(��X���Y�L�O�BD����n�Ѝ��\vjG��xh���6�.Z��bQq*��?���!i06B�P&��Yv�����HmV�L ��m��/��|���ǉ���������e�J�έ{d�r&�8}9�}�}Y��~!�����l�0� �·���E8�aVBv6����Y.�� �	T���0�t=�����Eb�����\.#�nGm5�\U � ����e�x4C���D�(Eˇ��=�Dg���-VMv ?`s' ��TЗ�`(W��&��_O�WDӾ����N5o�\J�W̨�W"X����^n����-}�}s�N�	���X5y�A�)��[��Z]P�)&sW���J�:Ao���)�#\ŅZ�A<l�sگ���Q0Dǫn��c��s�W��j��/��?l)�y�������anU@xc�����e�PW�V+�{=���Ų�l�H(�b���OZ�UϏQ��a}0B&gO�Ib�bT��Y�oE��P`�#cQ��M
�z��W��V$d�݁DU�Gb���vxȔM�M��A������=�\��R��	m�ۧ���M8&0;�)�A��Y'Q�S���cbb��v��:�>)�쇠[�FiL�T��0?J�H���e+��e��,�1܆�7�vݐ4�Y��;�Q0֚}����Ym�**�0�Գc��ԔY/b���!Z�w]}���4s
k���n��'�L4�w�BT8�'2aƤ���l�Go;�q�`^X��s�����D+񿇡(���
��ZN�v����z�^�m���!@�b5.��W�w�m☱��ڰ�c�V�(ޔ�W+������i�ǩ��d�3����>̡�Ʈ��}�������J�Em8���Ѻ��[P����l��i�>B�Z�&u]Zy��r��;<�xà�
���oH�%��>��9�)�&�*��m{�{��Efp���������5�����*u{ H�����>~���D��Q1��x�Ͷd�u����u9�!�A�G�����*�Ҋ�K��/����DNL'S#Â��SS�
��}ĩ����,(#h9	�ߡ���:�<�������
0�T�!Rg��C���@���A���:�y�:ss�M<�`�d����D�Q��#=Zy�,?޼ T1�wI����|D?��$���<�j�;7���7[�x�KUm�)�c҆\@k�j�wG�=���t����ff�����ɺ�1�2k�1jF|�pn������;>u�q�C��h%��;�������x������į�:�aē�%�����q/�tXȓ4f�z40��|9S��i�D �i���I3n�l�G'�+9`��喝�|,>���� ����`l��wQ����$ҀdUtLU�w7���ԕ�Cy��Ri��t�d�5��9z�nh��(l�O�K���)b&��[�hG3}���p���+�mO#���|���Z��3e�CT�fi~��|���{]`�M��d}B�㪲{�
D~�P��,��O��6 �&3(�#�A|�ؓP�-[���6�4$"�&ѭЇ����M
�&�e�)v���Boǫ����S�jf�X|S1�vG�kt�7(�V�Q�7} wyǰ��r_��6�Z�X��c��Z�i?n�_�uQ���5j��\��&�0�6Z�گ<��ޫʬ��5�9ӂjwH�Z���J9�I;��є �'~�o��b:ϟ��kk�|ǵdm�bvb0���sд>����-��'}ٔ��S���n�G߼B
�����JϥD�����8ys��H{�C(LĀBX)
����ږk~��"������im%��3��Q�E��.jz9��P痽L�?�:!�X����'����=���ѣ���{���6-m ���51J�Y돈q�7��\�b}���Ɔ�i�i�N�Xi\&��6��P���is��P.�u^<䆛?�
2�/�^��D%���:NjQ�Uh�P	:��W�����>�; �kK[��ҁ��#��
���,��SI	�Xq�KR��Z=X߂��7�{Or:����_�}�b�BQ�ž~�������/��� )�����^Pĕ7E5�i�w��;>0_��@B��
C������A~�.W6Ⱥ.����U��u_�{�V�Hى��]@�(���� n��4�8
	XnW�p�����)E��
������ߋ����#��Yg3�*v�L�X�#4�������b��Z�˾��΋�gl�#�蟾5;a\��j�̥`�$ڊx�j�վo�'��F�5��0S�����(#��ca*�&�����LV�t˦��Ĕ����d�8�nS-� '�4�X����]U��>Ї��D���6��=�j��6Q#>ݲ,��Pu=���d��HŌc~W�x��Al�7��6@��p��^+Q�d��7��CJMbJ g�41�j7Z$(U��/'ȭ%�*��&J>T!?ڥ���N�E���8A�� [%q ����'�9-d��W<�=�ZԆ���@�k6�в}�^�G�b�7���MFE�� ��q�:~��X��3�O�
�O��n�-p�l����6�i��?a��*|�����7���M:��7�z���l_�J-$$)��;��!�	�i�</���$�/�⸰5;�D��»b�&Ӣ'�E?1:�fC;�y!���_�JG�����Č&<�yd�(���w������Δ�VҠl���B9��T�=�Ʉ\tzr�E~p�ue���{Ni��U?�R���IφY޼�U"�.�a���� ��Ї��\�5%��i�l|�5K��Uͩ���mkg�lI�l���$N���ʭ�mS����lN����D��{��\�A9ïv���w��$��_@﨨$���ǌ�m��q�
�g�Q%)N�9�$�������g�9uCU�u�Q���	ʿ6�>�:$4a�,�5���ͧ���$���*i}W��C�n��/"��Q?vKJ{������6��;w�p�+��v"�7{�������-�,R�+7��{?��<��w��@���,G)�XA�4��*�ޝ�pd3��eŀ����j��M���|�<�c���n*��vV.��1�׊�YA&��b�[���B}X�*�'z���kF�Ȏ}+E�;���K��;b���\Q{G S8eǍ�C�b�Է>�W��$S(M�t�'�b�j1+>���;1{)����^N�V��E[�m��O��Q$T��+@TJ�M�J���R���Mκ�yA�l�45��)p�W+'��9u�u����+�,+۹5�WX*�3@s���������]����$D�':�GD�GO�`�`9��z���,NUxA�� ��G�&��Sy"�-���n��g���r&8b�\Aρ%D����&2U��V��mA���������O��]�R�d�t킀��w���MӵI=i�x#I���&.��1�UbxO[G��Y[R̗*��M�6����F�&]qX�o�˔MS�feC��;&�����Am�
��}��҂Xc����L��:��~�p_i(� N�N�z�(	�,] R�����i�]t��ZFy�;��1�F���$�C襅�^P��������H��"��A�J61�3t>o<�*O$Rܲ�B;d.b�z�F��-�y@T·���C�h��TE�	^�Q0�[���[Ͳ �7?��
�L�������a
�r�iّ�"A�c�G�U�/H铭���Bj%�m��ނA2�	׮�ƌ���<Z��Ֆh��~O)#&��B�0�3MbV^r~c>8EIq@'� b�6P�Nk��z�r��w�����m�����q�7p���rW��$����k+՗���Zʱ�4�9o�����s�pN���x�N�ur@��w��Y12�ҵ������a�C:Z�g旴W�𳤳>B��>�Nv�b�K�^8>�S�$\�H�}xM6�Y���k*���~�\젎�~��|�+V������;��P�,�K�"=�@r�3�ޝ�P����z���|;��F]��ؽ-x �8�+.�pD4|W�q�2�~�ÜH�����}��v�b6���~�d��E�_dB	qI-��(^���X�HF� -�̻g����^O`�f4q�����j��6��k��s�g����0��z1ą����ǂ���t������!�����P��;Os�Ui�BaWG��h"#���Z_ڈQ�`���*���f^�J�ɬ~���c� �A�F��#7�k;���a�+�%�����ٍ�(;�^}~�E��1㛽R�`#�n�U�}��KcF��Iz_D�D�;ttSG>���������Kb��i�����	��J����Ҕ
����5"
O�&