XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����0�%�2Q��yѿ	_Pi��3�l�=��ѐjAw�K3.nR�;��q5�K]]���Ah��U�H��H,}��wjV�7�Z��L��Tw!಴�ё 	:��»�6H�����[_7Zxr{�:w���	Ic��H�'u�j5�7��e�mR�g���W�;�n�����"	�Z���N�V{y�2�����˦jX���4���,/�Q��hǯ�p):Y�5r�&l�=tAl�#�t=}��8��6�%ߓ��ٲ�2w$�s�_�
��9����ﵣ�aIϮd<�̷�cp�!���ٱq�9tTy1�ZM��j���ǜ0�7Z����N4�{�0���|p���"�@������Cߡ��`��JH��9�r
���:}0W6W"�:mqZ'�k�$Ҫ�_6�Z;8PD���ч���6�b�.��W� Uc��L/���fy���Ý�d��;Z�>�{���G&�[�To¾3�p ���ة<�H�gNˍ���kXf8l���R#CSȜd���2m_��� �́�h�f�.?�c����}q+��b1ǣ�'58����N��͚�Ƿ���P��I"�zPf&����$i�!q|%vV�L!�Z�Z����<� A�)A������`�,u��x��CQ'�O���*l�ޗg<�I�e�G₫�bR8�u�mr�����\��P�~�8���ץ����Q��e�Sx��>|����ڇٛ��F�AJ�L%A�Y*M�{W��4�HW'afn�Yy�mXlxVHYEB    1d59     8c0%>���;n��4��-���a��bIB��%Ar�Hࠦ:�ը$PB�%��h�JA]a0�v`�O�n�Ӥ�t>;Ҵ~'/F�x7|��´��-Y7�E�����ٯ�A�b���d��t ^�O��`�@P����y�@�Xl4�/����10Y�͡��3}*m}�iW-L�~L�/l1�ں_��J0��=(�d�H	ʭ�i���V���P�Z��A�!��ٕk�5�~�#sM�R�/>�� �F5SxkV�ΐ;GT�N�to���m;�"G�oOrJl�g�c�i��4 Ě���y#�0|]���B�	-�'Y'~��e�s�eZ�W��kD��7~OX����;�ܬ��L	p�Yp>�2��6�sjTG�>'61�d�
4l�9���Y��&�!`���G�d�F"nx�u���qEM�\�5��;�>ϱ���8_�����vڤ�.�T}���퓌B2��,����_��ڜ�>�1ᢦ\�ya"�}F,&nI*>BQ}ۺ��^:���V.>�3V�#m.�)�O��s-}fЁߋ��JMU�j����ܒ��a�6�
�I>���mn��`lř�����@'��U?(���4�dD�F�{�+ZA�ˁ�A����|�0�I��	h�{��c�^4�÷Ŵ�:8��L��	_OI���
��h�u��� ya����o_�1ck�[���+P���	�Q�$��lb�<�
0�;k� m�dt�@�F�x�	SE�B���Q���+�(��Hb鋲jI%�y
�͵��7���;X)`��A���M$����T�n�2�%I��� ֋ć��?m&����x!N�A}��O
�4w'/y��_�z7�,�JA�f�Z�O�G�T���vj��q�֏��`��7c�-�,k��x԰�[��b�+rѩw��H����+,�l��,)�'���3T��k�8���6�\r�BL@�:Uij��CN�P�?J���z��R�HպxF#3�N�s�;���
�(Po����ub62�5�rS�@�'��M�����5���N���^���!������1�S��1[������>f�+DEtW&V�rЃ��f�EP�O<�I�$��y��d+����KB��W���ʪ{;&�u�);�bn�T+��[�r�uA�%����Hh���>V/���(�v�m�eN\]f��f��K�xs��\Zf��g�:�=Z���^�P�F��1B>������y�;�r\P��[MjD��(o"\r���0�x�8�X\��#�	��;$R����J��e����^�H�9D|����a�^A����k��[ɻ��ʖ�cr�?S���w6 �?DtMf�Gm�2s���|6��@�ZIr�ҩ��s�:�xl3���,XÈ�H�\��Q����5�E�;A;E	x�,�� &�6G�Tc@��{É:���:���^/�����D33]s0�Z�4���4��T8�z�7���n^�Z�͖/��Dtą`��P�X�ܟ�<Ȭm�:��ދ�Y��s�9����H�:����J�r�p'#~2����p6�$�EWp�%��a���g�j��	G�^E��������مd�j6��A<�I�<�|ɴ
&�h�0"x7�@�F��
�_�����&��^Y��O[�/���ݥ'GNn��8��e����.
��~�q�X�~�f�ٔZ?0d�ڏ��}�D�bH�pq�ym6y��X>�W&��M2Χ��Fu�AO��ZL�]�` �E�7"kY-z�b��Hhx�>���$�����pl<��:�W �<R-��pTq��8'��S*���N�������`������rJ��+(��V��t@C��q���p���Nl��G@�	�W*<Z��x
�j��#��Q�,߮D�E�&�2�)ȣ�u����C��)�*)\W�Y���k�9Ǐ[���kV�L�^���KU�8 ��Nސ��+_s��.r��aZ�"�o�dW�g��\�=膓��k ����s(�7D�>�a��lWb�({jXɚ  �.�Hi�vU�Q!����{��X4sN=kB ��h	2�W95"��C~#��U���0���z@����\ZL�S�&_L�/.�
G�4+�S����a#�n�r�@JW�H�7j�qE���K�௽�o�X<�jD�iZ�WU�8�vʧ�5���`Z���f	/�����*�/uV<dN-I����m:镞+θ$���G�������=s��`
��.