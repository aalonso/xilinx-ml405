XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$��A��@�UT"�NAL�6V��ƍ�k�_�oo�JI�Z��Z��K
����9��V��t,�_L7}D�c�C���.���6�Lc�3R)KBN~���)�t�Z�';:#�1L�mT� �*n�)o*�#!o��m�~�ߣr�Ң)�ـ�=��4����@�����&���
���B�$/�L��Hh7т��Q�1��{���}��� 9jn,T]R���B�~%�-��Ov�;�M3��`y�P��}�`X�<ÊpofzK��x�V ��9. -����t��c)�ְ�o�[`��	�庄�JXԅ�l>����0y:���YK�li �#�{��ؕ.eE�wl�K�;e� E�Dd)`tu���'�]�_X�E��#)D�ʹ��C��'�ȥ�_�l����`���`��<%�!�r��"�mpô7�4�Y��V5|U�A̮�?.�û�
n�g� /21C¬r�h �д�wf.�I}t��v0{h�6^UA�P>��|}Z�쇾��X;��ݗ@�Y�`���X`w����j���
0]�w�R����8�� ��aZL���K�"�����Н,���$��W�&Oq�� �bE�bT>L��O47�석<ik��
)��I2s�����*�B�_��_Vf�.LǺ(��#Ь��u���
x	��xxH�BG+'��]@��e�t�35���$9�i�vj�2,��r�v�󞪏E�y9t(���DW%P/�{qJ����>\��T(g�@��`��N�^B��ᴸ�AXlxVHYEB    1001     6c0�v'�Ø���{�PRz��-O>����R4��^���rjЇ��w���9�1�mXT��-/�?�l�����Z}h���"G���6jW:�'�N���;q���*��eaTU��r�Q�!f�
���H�	�pS�Z�Ko�S��:�<t���ҷ��t��F5�L�D��J���]Na�k$yB�0U�	��W&�u�ls楶���>zK�W�"
h�QPz]���T�45�ݕǋ���\�7�4�apk)d�����g���"4ϖ��.,��?�6V2�0��EW��Ji7ݿ6
t��1��0�)7��GI�)�clֵQP�||�vHL'�=Z�6�����J�Jk$��*G�C}!��;ϖF_:���"�1�ix;F��B��/�u��%�F2K����?J�0��El�(�dJ� �O;�$�D����i�`�Y���f���H�S��Ԏ�'֍-D�@89k���W�=�	�[�D��x<%.�/oҊh?|�T���O蹮�e^�3t*{������JY����З�cu��Z��Q,�F �"C+��{v�%Я���n$v����O�1����BWC�1o��T�U�Q���	�D_|�O��T��pEs��c?���]P�GY�wʊ���a*�=Y�Y��Ae�qV���IDXa�Q��}=�X��=e��r�/xi����t���8%��c�9�3��2�F%���=''��C�E9��R汁�����Ԩ����x&�qR~T�%+������Jz��̿rW~�~D��ȩ��b:J�J~�ԗ��!�g��-��6(F�'7�<�yJ=�Yz8�KT3�U���I��+�_d�}~D}2�����k�1�U����/�k_td/����e��}=4uPq������4�W �E ��sRNJ
���k(�x���� ���jp�o��,�V@�ڡ���4z��f��XD�	L�^�wR.�iEfoT���;:��T*
k"�]@����|AU���֬~�k�ld�N|�2���AФ�(�^�]���9�C�9��(JI�j��B謡Ad�È�Y"��[�Gd�P��K�{��Ւ���,��[�w}d磓o{*	��@ف�u&����	)�t��*�Yeb:�8�l\��(�F����p���yl�}R���2b�UJ얱'1��,*`�=�cj��m!O������/"tӮ!m������O,P�1�ڞ���K�<g����S�z4��W�%�tl�@�	����D��>O@��s"��WQ:��[ ��{Z�n����Ⱦz�C�߬"����e`Ď�5�)�i���;���F��0�A4��dp��^�c�~��w��e��9�!���&Q�𨄲:����z�7ˆ8+���c���!g�A�3l
QE3���V�Q�� �"�n��x�،�g>8�����mo�U7����p������Ai��:�jNU�o�1p�w(;����u.�F "��=��?A#��C��Keعh�T��Ӈ�|�-��t[���JC��\<	Z he�@���n2L��e�%M%7[�Q+���������^cJ3�Py A�5�Ss$�oA��}9�~�$�֑����b�ɘ���V�^�����]�<������>�L1�?��Af�h<�Eo|=C�%6�����}07�E����~�A6���J�	���g{o�efUشOU8���J��r�/#���7��]