XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�{
��e����/s��M�����r��ƴ��vk�Aɮp����X6� k��k��a��n����-Q��)|�5�(sr��@I���K� ��Y��Y�Y�C��a�]����_Yp��ǭ-�������F��nȷ��Z�����XE8��IS*?�3���9����{���9e{�)�2��9�紹�L�p�hm
C��&\��Xu*�|~��Q�8*M�H?��;~ा�(�'?�[�����3�s��`2b)�����$�D��j�Hlq5�����+>^|�4�����|����6{K���G�>�!�TM�kڐP����a�>��&�#I9��g+���﮲rт��/�����fa_]q��W5�@��������|��#�S�$��b�ξG�_ +�c�|X#�5���%�4�7�+�6
��%��֫
,}ِ���8K#�9�{��\��s��'L��u���O����H�����1��Y'��g0��+�0Բ;������y�[��<�/��֤M�ol"��~�y{�0�q�������}��V�
����}HJ1�)[�߿�s�ɜ��5��t�|=;蘘��X�{� 1<,���_�ǣ�֋��-6�.�ՉP�򙪨W�қ���K@�!|�Nj�����c�� ����W@�'a�-vq��@�/��8��Ē[g%�0f��L��6 ��᛾�, ���}}�8�y��|�8�s���ӫ=W����o���{����x�>�ԁ��tXlxVHYEB    4548    10a0�#�e���cb��^��l#ݬ�������h ]u	�X�����$�����[;�������]9�6_�_��xCﱅ"�ﺘ0}�:��Fn��2��~u�ߠ8r��6���4UFV���g076���?N2�&�J��?u��̜��a�ћ-�⽄_0yp5钀�N�@��>ƤC��Gh����#
�J:�nH����P	�)������p~*FfW��h��bl�Y�-�������K�p,�_�U�e��P��&u��s�渵 �ۯ^�ncH�r��:j�AX���x�	�ڹ�i��X��s-����òan](���GjY���@Lz��`_B$D����H(+��[��(�������2G������GԮP#0�@y�EH��䌥����Nhu�Ļ�$��Kc�dV}-i���;�?�(O�nB0�8�����m�M�(}����!�	�"cѽ�S��P�����^�'5t㏋o�HLI���#��׮K��.�~?*�eNv߅�ɠj49-�M�I��t�/4�]�!n�������'{2��u)|�~�y�$��Ym�F��`	|Ϝy�3�BԿ�u$��M��υ�
� ' ��{/}CAo^/�����M�wG�bs�8Y,�*�A�R�D�
c�����f���� ��W(��8�׆�Rd��?���ͰO�Y��ȁ�zR�з�����Tc�|Z3�{ή�� �zR��	۷� �M|yJ8�N���m�s�`�Y<��ӈyIeR�,Ct������b9�Ed((�h#�e,���3�}H9XO���5T5���v3��r!�/5��l��>��l"���4\��;�2S��]D�rm�:�����D*" l��?��&"�E�Q�~����ε�˓�Y�t�d�n���.�T�J7�_�7g_:�l�����!8�XȰ<�O7w�M^/��L�1ॄ�ON{���0���Ngљ��n���+O��F���a����'���o���%L+��ᖊA32V[7��^]38���l�׼�~����<jb�xg��:��wr�{=}�!��S	^��Xq�}ŷ+MN��D��s�2誇�����@ 7d*��.�a}W|���Z�n���ۼ���@r���{����l�H���-�Z��.����X�d����0��@����|�OC_�����t�^&.���=d�煅�5�d�Lį�UnK�A�+�Z�b�@�c����snL�,��6e%�\�lw�����1����U�2��c=�?>,o]qx �+
���q��WѪW�:0�*��3܏�J�V�<�#�
�	��3�8�H�������偧�=�Y�k��v��S w����d�x�>/��z�̵V`�OP��?�or~�?fpqJ�zw���
(N I�А!%�.>*���jN
,��I�f��)ؔ\R��@�7��FկD�3�D�P<��i^���m;mV���N���\����3�X��5�,�\��~R&� 8��������.(|h�N�ۼF=�c �>����炛���]|2�.�Q�"`��t^*�0MB)��Lѣ�ü�M\Ue0X� �h�d�x+�7��\[�?Y�����`�k ��@��KS�K����07�.Hֈ$���&@qt��}4�B>��Gw��d�ҡ��{󛧻|�)���4v�T�����ٶ�BH��З��Ч�p?A�����X�Lhd�o&ɝ��5֍�H�\u�8�/X��</��̹orL(K#c���k=�j�;��f$�ӥ�Ӫ%F���D[m��}�Hz[�8O�t���kH ��g�l�[f�"F����m%Մ0��2P��g$�Z���}�@g?/!�N���V�}�x�f�G����KGɌ� �� �
��b�U�TZD62"&���pqzO�ޯ�ae��wQa;����bĒ�k�:B����������4˓ߦW�����=%�+m{���Ks�}�@c�1�aڅn�\��@�iɇ���+E�4I�Ԙ�<&;7uφ�^=_�۝���G��`����늕��1�a|����O�	2�!PD7��r��fI����Ew�.Mu�u�vR�������Q�?�^B���0<VM^&��#�?"uX0�v�f�|4�H����y�1g���:�w�٠x ������9C�R�qxq}`���� M��5|K�� Sp��Yp@G�ҔJ�����~���[����u���J�8=UP�W��c���M��:r"��A$�#�E3w��ZɆ<��i�2$��k*rܧn=�O^.�K���j�.\�H;Ⱦ�$�k����d���t{]N�4���*k]�n*fs�WA�`]#��UĄ�����ԗVY@����q\�:d�s��
�Wd(��v̊���}j:�}�-+�6f�4�����vQ����瓢ˏf�o�o��z��N"C��@A�ߨ+!\�`Pw�>��\n��>gd������U��$��Q�74��Oˠ�H�z�u��wA�����顩;e�U��b�D,鸗٪
�@�A(h�D�L�ya*Kf%3�U*�*�SD�d��dEg3T��,G����(�$:��pv gZڄR��tk��7��F��놇3e���~&W|�^���i?��}��D@`O'Ɩ�gR��=��q�6v��so��?X^L�I�Z$����V�2��l�9[W�������+�n������L�J"����\k��k�^���	*�<����U/�LP�@�R�mm]ߟYe���x�2�tLs*��8dS������u GimF�v���6ŭJV��[#D{�j��J7@>5�qU�|���@����	#)-ְ<����p>Q�����[7O�AuӃ6g+�����M@�''5v7��V1�K�.�*��tU:]�Z������v��|�HJ��Æ�B���W_&����}�،Yt��S%,�����&��Ns����4�T���a˦��.`��&��o��]��:�h* |U%�uw�A��Ģc0X*!�ɑ �w����O� ��j���W&`�z��is���z��<�e����V�̂0$0�)����0�!)���`��DI�uUq�.1�Yl�b��lw�}W��HK�즻����٦��p!0S�� x @�tO��c���jXv�N?yt��B�2l�LǞ��������j5Fk�"OJa�.��L[�h�OL�_���$��y�~��VX��2ʽ�nX(R};=}�I\�wJ�X��T��!��ѷ�_}d��d�N��\</�!F�/���&�A���Dq|5֙��ͨUuL�>�,z�4�����s�2O�12�I��{J�#�����a�"tN5������k=�t��10/Bݯ��$�ů6��&R���`�ٷ���z������3(��(�:���2�T��]�S�J��ᒛÈTjEj��(��	��� q' U�}����a������8B3߿��t��<�qD�m�ǁoo�'���˽���V���6����R=(�/�+ܲ
������=�.֯Htp`{����D���TPMCD-w7��<�tAis���G㰡�QQ-���_8�2���b&����z> �r����?ؿ�Ͻޮ}[����>�k֝���B���鄶*�`��4�A$q�c�xwߝ�q[��
��۽/�1C�:Id��9���Q�Dx+Կ�L_����y-�X�~��I20����?��ܢ���Uf5�����պ�	$���$�E��zuB�o�����F�B���4v�+�Ã��}!$��1��c��\%u�1ĵ9��O.�n2�Q �[��-T
c�_C�o�Q�hh�@�X��{�G���\�<H�-D���}��hF��>f����ꥥ��c�`�f��!�$�o����p�~���.�Nf�;����h'��i�g�pb����y@Ú7�� ��CK��>���Ȟ��b��-����L#-+ av.��]&��	���3��{��ɢ��Ҵ}�(�����i������|�:+�>�$jm1�6q�BB�b�QN�<�r��"wO�sDdO�@�P%0u�u;��J���4(���Ec�8�.#�Z�<�|j]���A��z�8'S�Q`s�������ë�e=�d�%Y���Ux�q�;Sߩ� �����1�?/���>m����A!�;������\�殧ߏ\�QP�Q���{