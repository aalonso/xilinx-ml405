XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��՘�� �h�i@��l�Υqg�����({ė���z� �_�$���:=� u�L���(�����lU�S]��nC�!��&�ecC�q�Q�Z^�O�T�8��l��<pVA�bw�������$m�/'��H�G��5�L�J{%!�vk��a�s�Q��2k�SO4�F��8�Yw�)}���_g��V���6��k�`,lJuŭ,���wn%�>��о��Z�^�Z&�E%M���馲�m��5��PI�x�=�>0K_� `�0P�h)3W��wAz�o�A7�������2Pc��S�>�������.�Rѧ�I=E���g��.�S�KL���%lی��h�~^sS³;	�AQ/�^��+�
�"2��ŀ3�T�I����f2b�d���=���-��Y����n-���1���~�*�S�j��]��H�K#C�}���vG	T6�(��@���$Ѯ�!���$5�Ӂ�0B����H�Df���c;/��V����J05��A|l̽g����Q�M�,ў�D�"����顿������$�9�97���A}O�:�a�T�ƥ药Y�c��4��wlJ�i�<D ���t�F�!��<D\ �1�y\���@�4H�����cq���{N{���չb8�'�ZY���A7qaL�F�A�Q/�[Ⱥ��3��dT��C�*�ge�1�ӁF�r"�4�;)aK�C��г|6�a�P{ftNWJ��z+�t2�D}��݁{
�4�����L�m�:�_\ZGM~�jXlxVHYEB    159e     7e0�V-]�c8�8����k�"�G�m���*��cY�N&GP谔���뷍	Ǚ����DN�ԯ�2�Ɩ0m��I��޼C2��%�#�*d��"�Cq+Zk�����.�wG��E�Y�T���݊ [�Lk>�}�x�	�w"��E�1,��lO	��r_�<�k�|f�3%g�;P�sh~�3`g^��'� 2��T>���ů��e/~��jh�n����x��y<;�]���8��lC�6C��g�'��@x��/�M��tv׌S0B�Z�.K�ܭQu�<����W���e?�ʸ���m��PTۘ�\����`3[a��,��v�����&j{��ǭ3\���3+����W����+bc^b}��P�xHE��H�:�2L|4>�pXַ(�R"?�N$��{9Om4��WBhuV,�e�qV��z��P��!�C�DJ�u��^W\�T�6�Cm��0M釩�d+���|%Zsd��{RX1�s�V���a��K�h9����sv[������#����8b?dR�|�9��x4Ф&d��_�cRݬq���3B��]��C2Y����4p��c�T	�d��RNt�NnFG�yzQ ��zT�yigwD6�CSz����i�ލ`?�f�y�<��7����FGN^���u'��`���y�Q��I�sv����Λ�"ï�u7t�ڐ��W��gV��a2�'A�B��Jdh!� ��QppoM��1/f���O�љ�އ���L�ӎ�V�Ψ�gyNW�4hshNQ3��M�������\�`�V�t�t˄p��A���V6�oS�:j&u:��
Jy�q��fb��*
�7uj/ntG�_�C��a>�|>�qjɈ�i$���0��8�|*o�w������`}���e����x��R��mR�履A�$f�=�9Ӡb�����yly����ɚ�]�(�͈FG� ������ �Py���V_��If�̘O���zU|�������¤�ѻ�*�[�0�1��ʳ
 I[����@�6�x�j�����J#4�9L�WPp��q�1�Πsy	��1)��ux��K�|�+\�E<%y�TKZկ=�s!�i�|�M��h�`m_�܀nY�T*������g��ú���3���~�����1�+����2��`��ߡ������- D�S�|߮)r�З�|�D
P./�I������w�uO�8Z�dj7�����2�K�?)�l�f�p�,���ZqC-�w2��v �Π�Wʖ/D�<�m�a�p�'/Ĝ;��[�|KP�H�<0����;����@�{��c�#��̴���u���cȅ8u~\���h<��}'��1�sF'w��6��Zlt��.��q��\&)z�U�92g*3@���k�Llddi ���N%!��	����Ě��a�vc~f�s�TI��V���̓ފ�x�V�%}�g2v(B��8����������B��}�(~��Ѽ�|s���Oڇ�������,qn�'�Pʗjz�u\�Nŧ�tu0EJ�|Qى��(���j��:��o��C.`�TKtT�.��Y��%N2�Tm/����E�@*�ګ��Sp'=�>�!ޗaI*���VZ�4v����]�
h�?&û�ӪK���ĳQ�ADGlO44�A{�bݖ�Z��哧����M�9��V��w8���:�5L�=�<">}�[�	�S�IѮ�B��H��ǹ
H����j�ɾ܋�omuC����霞�M�Ô��X1+��\�_��ί_;Nx�1�B��\���w|����]�k˓*�G'j���p�T��{F 礳PB�����cg�b����{���\��X���1 �_i�%�L�uC�)��w{���?RhLY����C̴f;�Y���AT���}D֠�~���Ud0�l�j�	��;WZ�+I	u� efm�����Y_��.�Q