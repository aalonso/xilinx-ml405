XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���{��8^��o�s@�&H�o�>�{oP0���-[;���O��z9X��;���@����-�+�V��ڲ4<�PN�c<�"Ά��Y�9�]I��ܘ&K������*�O�����v�Iz�_)i����a�'�y�(`J�Fxd�`C���f���?�<=.U��}dSs�;-� CZ��lȭhe_��Sz8��ߑT��=[}��+����.7bc~v��Z �"c�X�6ue ��Y�<.�4@ƚl %Lp���k��AG��є[�!�}�x#e-w�K�,0��p#8�B��;h���m�'�خ�� �^ �-*;F&��+��#�rk����϶��~]6W�aT 5Rk����\5��*��H!��@f �̟I���p$]�_9�A��WX�a��,="�n��L����^������������-Lڈ��I�S��ٴ�P8{Ý��W�
n$!/-$/9����f�~(��Q����t'���(^��ѽ�N
9C����"�g�H���M\�OA�@L��+�d`�Uܿ�<�<_B��{�>��}Ik���QB v]���D^ M@rz�fu K\�8�+�pQj����d�V��z�̘�W�,�h�`��d��d�����|�����<�����vFR[LB��6����a�!#�؏����;��"��Bl�Bbg4Pސ�C���G4�G�1�� \�[0��b�>��q�8�(x'>3�����d�LřtF��T%GvpXlxVHYEB    7a7e    1af0Յ��@���9+	T�q�{$��!`���Om��s���39�3�3�:]�U�x�8R}���܌av����΄9}d�	&�C�DA�[-�,+����iK�A^�R[6�Yd���r���^�w	[Q��.���}ydF�#d5����̿SV�ʕ5���͡���k~hh���	_��?��AbE|B�p�]�$��q��{�ܫ�gOi�ԋl�G��6h����Ϻ�Rw�*�z�&CI��W�Xzq��|X�vJ�+i(_�TlX⃒P�C�%����Z�
F���0�*���R7�>���ө��S�*���'Fv o��W�&�P!��2������ꆚ�C�w��@=�Q�z���=M�x�Md�[�`�0�PY_�ۅ��{�Vb����R.��{ �W�`�<�ۘ56�AE`Q���*_�UuK��(?@�L���ˮ����'r�~p��SN�G�!�}E�Y����&���~��,�?}|�O-��2�8eq�h�ѩLy7W�H�+j�E�c���k��q�t4�_���*�<�ekx��)�dwp��1��պ��~l�1�[�Q����F"��\�0�'=t��'��,=�1�E����}H3���Fs�oM�~�
�yC�2�ޡ1���n/���P���5�\�Z'N�X��S�?u�3GɎA,i��+q�W���(�uFW�%]l2X7�����>-f'�]RO�D|�E�����R0��ያϴ�q��38�~�\o�ҡ�й3�Uy���{) w4l���x1�[�;}�~�i�0��K+��fja)�k������#i&��+��3?B���^�,7"���}���9?�O��F!(����3��ɱ��*Y	��F�4�I�N�7�M6�=˸|�l�����h�7vLڑ���f�a5u��>���^�u��5|�c���$�i��mn"�P�x�������zQ�"jg���5*��b�h��8��E��_SE烮
�a���4����҂��1���}ea���A��ń�rS3�8ќ)���hv��w�1av�3P=12%t��҇{��v�M������@���:|�`_I�x��&�:u�����&2�&RV��3K�mn]������0A��/�Pn�r(/�eJ5[:�o�:� �T=%�v��|t�s�&����=��"�oPG��'}���I�0Rj���e�8�|�'(��z��85K��;�%�ժ�~��3���UG�H�iRd1�@)>̷4���5��gqdc沣�1u�r]����
�R���Z�7 ��+��{[}F,��`��>a��g���`ү�������͙�����, ���yqPl���V"��'��ڝEa3Z񿛀}�ݦW�~_����;��Tw�=������).g��ά>^�B��ʿD�ѩ2F/I%��B���m��֝�
����*�+���̹z�-�ʘ�hi#���E��"4)���g���u<���<K1�|��`WjU2�p�Ϟ�F�0��4�X��p�����R}&�.��%����9O�4[�l�=��)��GQ��;���pJg��ӷ����G�%w���� ��
i�aĸo�j0�1���9'�@5"��jTI[|&4�a=��<��<z�����ܠ�a�j{He���+�`
��|���M\�u��A���O��/C[�h��G�w���tK�_
nX�cy�@�z!�R��=
���+E�&�q<�g��pIjA�U9s�!W|�-i}=��M��u~l)�i��|y���#RU2�Q�D�ݯl����@����GU3�m�%��,K�ۘ�����*Z��o^�[ف/��|��b�9([M��:s�W!ŗ 0i�.1�N�.NB�1�(��P��L�˕mX�q��Y�=�6޶e�!a� ����Mv1̏>P�'�{.�P�L��'_���w��7���̻O��;���u�+P6�oz�^)��ؼ�^DvV{c�s��`Ώm$>
�@+���S+n�s4��T�u&���;�rd�z/���m�q [�d��]�Cz
uD��B��)h��R�b�e����ݤ�U5�b�Q��I�?]Zf(/О��JV:�{X��33�Kr#<��0���`�hё��O��9�����f���@��J�L��{��3KĉL3�-�j�L�r�T���]eFi�ϋ�y�8�Ԕ ӄC�`.��]6/G]��װ#��U�ʋ��
��B���e��J����5��'��}��톤���m�ս��1��Q��Zζ\I5v����:�n�3\�+��΂ߖr���؋�p;��8P���8�������)  �Y^�WR�P�
x�S�y�\NbV���!?ES�8o7�`�d���q�L�� �N���r3�{�7I�2�v��鉶��U����@ʉ�>Q�DxՑ&F1U��V���ٚ1G�8��?�s͔��/�(�N5�fHh=>��9am�T��xO�X(�-�G�������~q��頕c��q�t?g�š�רN��(������u���G���c	�*��=���� OG�8S13�]�f%mv�,��bp��j7�;���V���'�Ԋr�i� A��/����X�P��xjb�Z��$&#�Y�ng�6s�@A��M�� ��'-��v� �m�6zBh�%��w:@]�A���뜝�	�p�5�5=���H�Q��gT�ؕ�,$0m�Z������G���CW��֧�XU�Vh��Zn<E��[b*�S��k&­Ϥ��lA������3䳡�l#�t)7��P��)�$�]F��H�������0H��sd�t+'��s&L/j�A�>�s����CGM�i�V�re�k�q�{c�Rۆˈig��Uk(u<\r�ik6�m����F\C����橈_ȧ1^�p�>���]���*�)���U��^���T��XF�s�)�����q��f�z'Xb����Y�-ko�����8�g5�I�o�j7���%Ĥ���f���-�H�T������ٝ!�ш$O�H��!�t,�~y
�Ф�,/�����F��7�tCf��=KC�W$�ƛN�E
Q=3+�˕�l�&O���;w�����ƿ�Ş,�|�U�u@�Uٿ#���kۼ���ڷ��x�%���9Uܣ��+Xg��B�� _�{X5b�������R����n/� [�Gs�lY�[!�cG�u��r��a*�
=�N(1ύ�[�V�,Ā�;�ٷ�dO�0d!�	�&��A��oT�5�B�9�7��r_M�{<�"��q2�y�wx���o���JT�(���@�����9�K�~I�Q�_��ۖ�v�%\��/�i�m�D�b2�@����]?;Ә���z	��SL�rbπ�n��}��R��0�j����J���F�:��_XW둾�8y�V�*{ޛ7�J��rEi�
"��f�dQ3@�ӷfu��Q�J���!� a��Gf�Jw�.܁�%�Q�6<�'����P��"4�{� �d�Q}�����=*��֮~e��囕�]�]m؟2P@��U`��"F��Ug����U���4�9�k�H��[�u{
P¾�ס��r��;�����a��s�G�7рR��X�*A:*M薂��\���J]5�Έ�U������8�)8�_(ڤ��_�
I.u��8�v	Y9� 	c}������#k�"���F��*���+E�4[��ռk�V�������{��9CU�[ۆQ�	��C��� tI#�1��w��t]Ő�0o��E��C�ܚ�b���K)����|�������̇���B�ǎ���f�'>�4|������v��g�7aͫ� zG��_��
G���g|b*5jV��u�ѝ�1J�R]_E�Sr���^�l�*�F��/_��������^al��KlGk�$��w�WLRb�3���bH)�>$5�?����R,�s�H�X݌������럺U����G��]v=��BI2�	��Л*��NK��x+_�I4%X��xds7�fU=�������y���N����.2፵��P+1e�,2�@�w�`����X%�H�� �J�3��]�mk�V�@1�y����K�r�43x[���2�����AmXʁ��͠ufx�����\�X�?�و�B"J��6딉��D?y7Q�3�آ��#P�]�t��3"%,Ã�
�R�-,��&������[^�\vn�5�iR ʥ?n�8YMC˛���.*9��R�||��p�K�$]Z��u�pwx���խa��Z���h�$I9���g՛�(�~�^��bνO�;(#/!� �o�-��"�?�1�Ч��'��"���I���[��N�I7ԧ?7n�(< ���	@�&��m����ʹ��{.M��x5�1��5���^;H�XRDB��D��dʾ,0����_�6�AۡF5kD�{~��Q�ڐ�Дr���$��p��Z)>mҝg�9��D�|�n�?����2�j�I�f��LL�Tq�ȫ�A���1��
_�S1�=Y�|,N��Z[��s�g����"�*I�3�$M���g�@R�i��QR7V��f�l�~]� �ua���q�t�賊߰-d�~6�=5�SEw�M�S�y��|��Z��3�����O�f f�WK\.���B�v{�8�ӕ��;՛�����z7��cOl��@�8}��F�3�5ٴ���Z�-�!	�Qd�2B�[��4����4��돰q�+����U�nd��=�$�R�v'H�+}󗆛�)ϙݯ>R�n5���s@e���sUOU�$�;M��_����W���	2Q�>�f�s�rx	m-Oo�\BU�!`�w^���w೗ ?�{:�.O�����bn����21O��h�l��9x@� w���z�2J����֠U��j�Y.6�<(,.��Yx%�v]y�]O�E��9�v��볘�c�*46]E�[;���yN��բ� ��c�Sw�n�g����h۟S*Y�D��?��u>l�g%�9�l���e3�No�񨱵Y@��Ur�a��K���Z+S���ȹ�} �t��s��B�'���1L�֩k��e�]��4A{������k���ȳ��>f"i� ����3�ģ�7Z=��e5?��ͿU���^�}���#�	�:�k�=~�t�u�4��b�S�{w{̕ߙ�]��Ǯ������V���}��׊���+͙������,@�%�V\���RP�OHm zDi�I
�Ks1&�Аbʎ�Uԩ۟�}�s\�k#!��y�d�1��r���"�h:]W�6��8�A3�ˏ�=R;!}¯�7���9��*¤��1_�"��ra]��Ӱ�F$�5�Լ��I"������WkYx����A����g�c>BE��w���%�~P�7�E����}�9`�G���A��P��y���"\@A4�^á���Q��/��2]tަcAsK/�Tj'٧�ܧ�ً��rV�Xe����2%���i5����Dd�U_弤�'�HԥL����JG����8>�Ye1���Qf���{��f�I�u��R�~�&E����W�{s�6�ؤ8�%�\+/¥I�6�+�u�P�&D�1��$��{�n�x�&7�MU�d��2�Z٣!Ӿؕ�iYvB��>�%��Ƨ7Mo���͠��F�1|�Yq���]�ŪV�>�&ҫz�Rl �Ot8B޴T�/P�qq�l!�u̷)���4�ў"�n���k�Z�+�ǌ�B�Հ@�\��� �3�j����o|�l����07�"�%8>L^bC�i���@'/xe�F��O!HG�X�.�pp�Yr�BUK��I��$�r��p|��V�����S��T����f�$�+�ş�o�m��v�$C}w=}�Q�"���`�;ݔMK��#��}�VQ�A�Gj$	�TB���t������V�v@
!
.?.߂���ȃ�וŚړ�i�/v���%�3	e�.BϺ��\�No��E8\��6(�Ho�E�.�e�}��D�RP�";�}��UͥL�T^����(�L��
s��%đq�scd��.�T�p���4hJ3��`z�s�u��:��B�%!��!��ZbR`�������.*�+=X����=�gb�,/I�:���9��X� S�O2�}Mxo#|��i�Qm	��X�_a�U54f;�k�'�@
2�i�M��MKH�- �3���%��#�������^9����q�U�?���Dr���9�RJe/a����8��q��7���l�ʀ�}W�5�&y|"�����5X����p�w@7W���7��dqP�	��Jp+���:�BK����/�W�m�4�;�9:߂8���:����0��E`+
���p~m>���ǉ�_�sYӆ1gd�D�xp��&�nI����	�,��)��v?��
���(<��ɶ)��j�C���'ݞrżF}g�rR0#d5|�X:��	J,�^���P�%�U���}P�z���;���1�/7��Ka��S�1Y�ѲD|~���;.�Ef'�<Y��	;���ϡ����{�v�]�����T���=O�*�Y������go-�%IVzǋ���@d�;�:������;l綀�UW-��=�±ק_����?w-.�5�F�я�N�gw���k�7&n4u%���U��_�(��{�4�K�(�q���	�E"��>�$$;���}�����{��N6�$�ÑH��-�'"���´��*� ��b�P�W�9�q�����\�����!3��ę��i�f�W