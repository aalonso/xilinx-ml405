XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��e��q��&��f�b �e��.��ӓz���3�se���ͮ��t4��1������σ��Om�<�
������נL�;�r���|��ͥ`�N_��r"�ȥ� �^�}m�O�6�!�&������H�Y}U�uf��`�l���yh`h��Q���5�nK����R�L1�7�!�dYE�N��xzw��ܯ�-Ns�g�%z��kA@j���! ��
���ĴCl��~$˶O0y*�A"�{MWԨM�ri5�(H{���L&h���f�t�frl��Ź�l�'j	m���ǁ�nutus�N�t�|%�Vǀu#ŵr�@K��1w6��!fL��Y���^�LV�SU7����/g↨��mIP�>��}�9��G9uj�wgZ-;�zg�l�ԃ�9Dd��[�T�	:C����;���#�,Y����A�.�#_⨦���=
���S�1Z���V�Wqc��
)J����&?��EaA�o��=�螽�nb$�B�����r5����c�fHɥ���>:��\[!S��SS�s$�ݕ%s�P�B#���*�36m8�S~���*�յ>��$~�m�����-_`��Ҋ6��$PQ� !�\_%�e&8��+�uV�W��6�<G�k�o q�.����$�~J�Uzn�e!��a47P��Sh�&�����`�v�\.L���T��{������8�5E"�=��5��%DbP�rwz?8u�9�U5�B��ټ��vxS�c�e�7���K}XlxVHYEB    203f     a60��X}m�:|�#��I�U�����zh&���4a��?V��U���	��g�/gDd+�v��m��Z?� �ǬB�n;p��yf#T�}Z�9�N+T&���',+;�YE8&���f�j�9�?�b�U6z�:�B������[�F��=�Z�ҍ�r^��������ԝ)j��D����9����W]��,�M���fe���[sԡ���C#�:��^��ͦnts��M�����gN&8��%�U�m��O���6-4p��s>���g-�S��H�.�	Et��${��W�q����R�5��t�"��H�6����J������Y�S�o��e��Ny�8V@��$�<��e�$�k˩�aVh���n{�y]��1�Nʦ��hUv�*A�6��G�'����|n`�p֨�_��t�B+V3��P��P��Ŧv�	�v��S�j��a���C���2<�[��j��~�G0)�=K��Y�7�K��d�V>���b�S&`J+ɵ�~�@�/��?�(#�Hn�]��ٳ����<����������B/�n�2�ݳ7v����H,W�11@1E������_����4K�jy
�]�.^N9����X���Z8��x�k�i���G��@��)�/�j��NHuN�K��&�I��h���xL&U���1[\Ē�́w�:�-�F�clv�5��0�ݦ��,f��`Q�v!��x�L������h�C���_�f7��CB�<"J��x�J%h�C=I��)`�C���w���?D�����#�:9܀F�A��Ra����ݩl�E�@�@8�q>�-뭧H�qo�Sʗ+v0�l��z��;�������|zy*C�����N�70;:ˋ�~�R��Nu��1��H�	C	���%���
���[�i�і���^��H��[k0k4�`�d�D-��^�"��2�P̚]�:����J�����K�0~%4��k2���y������)���dl��!�`��zg_*��kZ>�DFa�DJ�r���J��Ш0�ԣ8W��8�_e�G2%�5<�����kI��c��:�Ԗ�R�O���YA
��f�L��0�liu����l���5c��H͞���O��&7i�u1=V��MB�`Z<�*��߁���6e�L������/;L6����Ϯ>Bٛ��A�I;��삭MǏ|�1����S հL�Z��|i�������5�,�w-q��]>8�o�SL�?������9 �P�wMܕm�jHs�)c�S�m@Kdr=���#5����,���5a&�qF��ѷ�X��)�y��fܟv��W��R����(�ہ�q���;!YB�?O��HQ�WL�/�l&�+k��`=����5�������> LY}.���B����ķ�U~v&���RҪ��5��-l�/%}]�N���%��)MSr����+��u���}�~��U1��C&�����D-E�t�M���J�8Y)���j{� _�Z`uO�����@��r��-xTɌ���l0�[�LfI��[U�傅쵠�j����u������z��XK�_�̷�6.D%�7���bJ�D��T����� ��X�آ��j!�9w�cIv�N���
�o׎2R�y�͸Z��h��J�Ր<� �2k������^��7���i�|��=ۓFί��{� �ݰ���m�V��>-G;��$��	����=�-��E�L�(6���%G@o,u닟�V
�8ta\���3��%�)����@ ĀA�0-����Xyq�V�{<���Ct��g�\����&�	����p;�[ɦ�qct$t�$��y�(�-�]��u���T�=I+s�r2Ņ�1%1�6�7B$)�b}���,}n�)��۷����4���/�F=�'2W��é�Cz��xy�0^���<O�,����D�g(�`fqD��(���b��P�Ҽ�m:w|�v%�\ nqBs���u���Y[F��2(��ZW�v}�xLT�M�~;��o����v)-����"0�2�N�����h#g���jd��#��zx���-Z��i<�sVH�/]�p����#|�:������kC|>��ٰG[s�����	,�#,s�[Q���qj�FiZa;�.1���:�R�C��(�	�$��K����i�uoh���zIK)Q�W��B�	�}�f�j��3����[o����=��9#!Jj����Lp��R;�	-�KiB�$[�c��	٫����DF�����Y�"�3�2p�[�mO�^o鞜��_1"Q7д�b�v+toI~��xL|H��[]BI���lv�L�"=ᯔ>�b��hO��]~Z��T͞��_�-�fRK ����eb�U�e��ɹ�a�ҭL&$��g1~��a���,�sˣ��+���DD0��ϭ�WePq"v^�T�ԪE�g˓=hF|��n�Vj��7?Ӻ��`Pmt��%pUxTf*��lt��3=��f��>t,aEM0�|�V�r\/�c`
\����B�f�����Q�����\k��~|��K���9gY�L)���bz���ic�k̦{�1�nD�"=�o����1׻W[�P�q:���	"�:WAF*���p����mMۉy]�`� �����J�=]�[�H�&�	���t