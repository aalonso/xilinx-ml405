XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K��Wd�bq|�X�����՚䱘��{�K�bg�R��U�,����^�nO���O)�m?�ƙ�R�M��{a��J͔�ΪyiK�ݻk
n9������ɠ-�\��'�n���yT�-�����#9�U^W��p�x�۬+��IKu��M0;�N��}7�8]܌��;��:F�l
aɧn�ä�pϐ���[��N)�����oҎђi�]t�S	}im�����8ˊ췲Ɨ����ž���j��=}�{����O��/O����"+�����j�ju{J�+	X����$���g�C�J�7T��D0ϯ��u�[*�r:�|8����/�[��c�k�1=9�'$:��E��.u{h�'J��W���`ƭ��
��Kϱ���`� �_Y�f���!�l����*�1���PY����ը��x�N�Yӆ��Y��ז\0�fV몆�Uw��H{�:��B|:y�vڭu����X�	�)�z�e���"�m(T�~\v�4C��=�r-qhW������uGG��a��d��]�4XK����y
`��"����L��a=�c���5Q�= �� e0��j�R���J
����/���Y��L'E
�W	�	��35P?�<�`� [V����i�J0u�`�D]�U�Ȣ�����n����l� G�#���8���CꋶL�[����Y0k��8}��ks�O�p��HhG���
Y�c/'|�*�:�z�J�P�Ug�^~=���ܡ��b��cc`���\��	��w�XlxVHYEB    9653    1860����w`���� ��j�����P��L�YQ���Ƅ�щ0X;�?�ֲ��� ;K�nz��ul���8�M�Ͼ1#+b���p��B���[ k�����DM �\�\����R�����Age��L��ղ
����@|%�uu���ѓ��F��Oӝ0�xe��
��jF��;sh.z=��)�e*��������[NC�R�R��L�u����mA���
rňI�̿�z����t\��lT�X�˭n�!�J��m&�4�oh�)1�3D������>�%G�5��f�� ^� �X
Lb1	5 �1��_�[����ӌ���*e��J>��u�g��Xɔ��̘ND�<mW��W�j�-%4i�kl]��mU��.��k2k���s�o
�����Cw��v�ym���@�d	�N�Uy�S̻��TY���â��#=]��=ㅧ;i��w=���
OI����K�b^�0�y��Rb�j�OAIC�T�j݆vf�޷�{""><�Y35%B�KI��rc,pI�U2�ݻ�i�[���2���)�K���h��:�`�M�,U�8��D�Y�����J)
�un��*lG�^ ������r�Ň�)���Й!�>�W�A"�<�{S<"���W�
hOFK�!��h1�B�XIQX�tA���E���?�v9��kgԤ)W�'rE��Ħ����Q�ШL$3UN�{q�5wy'֧��t^��S����m ���YKf�˅pQ�WףM�h"!Q���ˈ����7o]������N�fO�����Q�wd!"X�[��YM�ɅE�D(���||��Y�,Śq�v�K�-�|��Q3�&��~\T�ܵ��Gr�K��~`�y0��X*8�C^��*��MW�~�֏P�&K��8>$1d#��Qb9˂�.�7�����;�-[M|��7bV��ڜ��y�ў���AY/�3�0�>Q�E,`d������:�H�<B@��7���[�j��;�%}�j,�A��M �XB��r�txT�Gܷ�P:/?���Γ��xw�prG'Ҏ��8�g��w�-%?��K����K���8�,0�����$Uh�S�N��Q��?͢y��4�Tp�H5b$ԏ�:/���'�� �3h'I��>�����sE���#J�8٢�73�B� ��%k9�NW��'���.ۄ	����z�Q���U�h�`�%�s�a�@�?&.�����c�^�^������l}��	QeIɇwy ��Ho副�V1�X/х�`�Gr�z;&)fY�*�v���I��5��g�}C�פ������}��^�X�/ZX�ۅv��y}0�B�r�������&�|�m� ��^��+�ʮ�
O��,Д����yד(�с������ �
`Ʃ�5�]TF��)�	q����z�܎w<�~؀�u������s�K�kw�ρ� wubD��U)dL�|�oєS��EKU#5�Z�	����ޡ
��<%o����{�m*h�˝�XQ��?C������)!:	��}=H���?kd<���I��RN��^؉�_�85b<���2�SQ ��a��X��[���U�5�"͂Ħ��t��{W2�dɱ����rZv�h�h��t,Ƅ�\N47ן�u��Ź�g���XoG��z8-SQ�g�s8����e�n�D[�q�>><�F,ұ~�%��z}�+�qj��!�⌱�����]��\~�B��h�)�R
mz���F����{� /3������Θ��@��3d���1�Z�t4�~�=��C��T$��+� x����@ 6��c��4"n�� �~rkv���/٨r"ϐP��ۭ�eД�[�]��`����b��<�X�vU�7�i�8I.�&�����e�{l�B���U"?��{��\�PvQ��ӕ��ff�ߡ�ꔃI ����4�/m�^�����b��D�P�"c2KciM���SB��;_��c����^=����y=ѭ���ߪqK.���梉�j���Tf��Z S�����\E=֏P�X�È�Ǟ��(W:�җq� �ZԜ0k.ދf'�`dV�D��o�ٵ�0�ą�Z�2���J����F�3
m��׶�E;t1:;��?"���v����:�@D���a?�Q\�=r�lWQ�(�7��j�M=�jUe��D�#=ĞR}s��4���I�m�[��A��n���f�>�P�G��7VvE��T�e#:��\�� ys߬v�-?ޠ��d4��K�����딃��G� ����,�a��QV�J	�H`��m�o)��'L��U�}�E���/G^�C'��`�0�ž��D��i!����{�IF}��i�b�}#��^��Bn�T��h�3����qR+�0���P�|2{�;��I�ĭ����;���V��n~$����Xݼ낷�1�yAq�u��rׄm �X{��+tu;��}2H�Z]Z�d�SB��o��{ '#cI$�+7�c�z�I�7_����;�mk�cv{[jЫzZ�v�[��JZ���q�
_)���דnLPZ	�
����a@BP�쨌 *��Wn�HvQە��s<�`�1N:�l�jJ�Z�X��|4όP��/n�40{�h_����'^�fE��|�^Z�lZ:8`OFH'$X�+-����������a��q˗�$W�����3�3���Lq��.�fౢ� _�gu9]q�R�C1h�M�s'S H �����㟟�R�RY���qᓉ�x��͉���vܷ{�k�ˑ˗h U��>��u����~{-�Q#�����>�o0���/���+г�iYr�н x� t�قXQ�l>�
xwm�wf���~+�,eM6T����^�U�S 1�2F���Θ�7�]�̖������y�>�AL5n|$��{0O��=�e�8X��p�S�x[����7�o��-��ܤl���c��0���n�!����1A�b��"��X�k1-��̀��aVs	Rt�Ղ���h^��9���;o���i򮱍a�t98��g���I�{�N�e�
��BO�rkT��6]N��ZJ�̊��k�-k]�����������
w��ZȔ� S�=� l�H���k~��Ț��揔�I�uJ��S�.��g�[7�Y��
�A������J^�jd�6����P73a�&��S�����
�K�c%�]K{��*�ӛ�"�%,82R"[������O��ש1
�4�6�v:�8-�p�~O�*�h�#���ޘ2�T2wO�q�T���4'H6HZH�qgQО��,�q��ђ���c�A7*+kYU�;.\�n�}n,VT�K��-��+t���#T�A~����eU\��r y]�*���p���ƬZR(��|8�Nڦo�䧼䰶X
��|u�Q�Ž�Nm����>�<�W�M��F����2�!w-a�k�7�T/�"��,�	Ѐ @�g��mOYbӓ��)zf%`;�{�LJ�sj& D2�>�F��%�.Ψ�s�c����%Tp�d�S2kB!e�vB�髠����u�$$վ󅤳��ՆtI!z���]Ѵ���`���}��r�y_I��Se����>�=��TU�DsCK-o�W��C�i9�i�Sg��^85ڹ#�;	�>;E ��a�^ycx'�C��I}���[,n�~۔D�d5��wY��Ui�D��JY�`�T�r�����V�zӻ�AQ��Z�?�^��~	�D-O'��'���U���|�^;6��(YY��d�b��'����o�ci�'%t�k��w�	mR]���a��N�w��"���g�Ldq��e(�p'��Oڊ$�6��^�;j�>�c]G�v:)V|��G���<ѧͥ��j���R��BWhm�s��C<�m4Q'f�ƭ xA��J/��R��?
\j���?�)�Ż'����۰��{̣��n"��;s�J�]���r�w���^
`֫"�F.MR���&q��Y�1��j0l����&��|���>zP��E}��|�(`%���xh|$�~ui	Ct׀�p�g���C0�A���59|�3:v��Cyu��n��d��q%��M9�y��i}S~�6�	Ĥ��#
4�4i�/�˥���Y�=/� ��l�׮]��UW�^`7���\j�t���(2��Q���%C�b{`�� 8��}]k@����}@�����J�[�w�*�Kw;5 ���0�Ȕ�Ќ�2�oe�?j̗��\6,f�%H��4�s�ժT���)����"���=i7�G4��:h�tG�<G+הbl��Jcc_4n�h7��6|�����X3���K[7�`>e��������cߊ��7�̚Y�8"b��%q�ڸ[X���3$���#E�8{^�ߵ���.���Qg[�bUm��p�/;�d��ʅ<�	2��bP6�V'���7�zwt�%�'�[Xtg��{�3L&S�t�3��$����=�ƽj6FA�*�7�=�2�����3���=��3��a������?��̓�W�$��j(���'�eE*���N{t�'
�h��Р��HK��r�q��$���uq)�j���}�X����0$+�F�N̈]�6�����2�4I*�wc+�R�i�jB K㶓��PV���GiAi���G'���e�������*�mK��*��3�I�����f��ˮ��	�"��i޶���r�$q� 9�le.�r�`�i|Î��]�%��#��֠�M��=Y�3�"zɞ}�)�ƅ��wY�8�,,|��TW��3����\����s�"l�B�/lU���~?h@� ��V�JKs5 ��|� �9 X�t�D�O���k��U4X�M��m��쉫����MD�L�ؔjEb�J\P�#'���E)a�g���d^���=�!yׂ*��\��	�:������K@��|���~� ����w���x��[�n�I���j(��yc���2���0�����}--�_,�Z�h�U�yH�8)k���D��x60�����#�D�}����,F�,p��zu�YF�:Ea���+q�������as�>Z�J�ֹ���<^�^!tv���}z��/2��2u�ҡ�Z��#s�-|�ʡ�@������nY��H/�x9�g�_^.�!�P��ň�5��7m<����X6?wW*xJJy�I���'��3`�7=2{�i`)@���zd;��;/Yn��gL*녝�m�� i�Rn�jԵ�i�	3�6�)����k#��!4D���9G�թ�ae�F4���f6�����W���3,j��٠M�4�E�����H߂�S�*SĚ��c�w�x�g����5Љ����X�Oׂ!�7�=�cE��#o�-���n�k}���e��w��32>�+��v�y�����;WY��C@{�����e��+Ҽ �j7�2b1l%;_�L��d]����cp��`I�du�|�NQ�ݷ
"D<�r��ŷ̖��,�G,�z���A�	R����d���5p��~��c�[&+�b@��
:��vb���骢sٲC̈́&jH��B�@D�{=�5��X�M?��̰۬^�ߥ\Z�6]k2�>�/��kt�[�y�����!�胆���9]�뚑{�=R]HX��ޓ<�MM�w����N�W�6ȭ���"ԩNNF����V��X��F|A8����͢�S�n��.�:�ygC��έ'�2�K�6-�S��[�/�+�5��5hoT<�Za�}��إG��@��dޚ�������|���˴��2.���ͱ�r8 Ua��k��
�EY���9��������*˘*.�]�s@Gʪ��}`1�{)���	t��Ϲ��%6b��p���,�`*B}���(V��|����}�;Qdh�,�`�ԎG-[6���8��ﬠӘr� ��+=��U��q�M~��q��nK�x�CYFջc�g�2���
���Ě^�_��Z|۬5����7�	[-_�"�}�iQDb}���8bQ3���Fͽԍ	2;|Ţ�ҠӢ����T�l�GO��)Ί��39����C:F���dϛl��>��KW����ܻ����`�ZQ��8t���O�F!���֥���w??����5j�� {� �G�Z�s(\2���,(����3A���