XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��O��p�rH�<��X�t�{�P�}?�itD{�Qz1�I�J��ǐv�
�a��晠���eL��뤕�ڇ��&Q-�*�t4A�F9���Ē��̵�n户.���\P���cEp�n#��B���}����	�����~`�=T�BɴTS��`d����.����گd�8����_V���8���5 �<��JH6K~eV����竁�I����L!3r�X7H�G⇃O^`�C�G*�:��o�e�z^H5����Y�:��t]*I�o<��/׸G�[�Z�I�7��!Pz�5�w	~8\���-)O�_��^s���(��^Z ��M\���v�d�4�
M@ݺ�P��/~���+�qa�q���#	dY�'}Q�C��cf�z�6>_N��1T��h�F5�8�x/�Nv�0��\p�i3�%��\��� ����o �V����1�o�� �T��|i.{g/fCD<�OwĻ����4µŭC���٥�f�R�~ƣo�^-�T>��E�qL�3�u#�!���8�BM@Vg��z'@�荰�����	K��p�1;-�*��wKu��ەy�m�1��������յ2���]�m92�J���%$���pǥ�v�����뼱�pW�K�N��J��?R�e���8��j�!LĠ
� d�0i�����f�$�����J���QxF�q�#�hܠ1 �t�v�l���@'�@�͐���'�=�!�eL�+������A�/0X�h_�ETd_����YCE8XlxVHYEB    5658    14e0�a�N��Z�&��Hr����[e"8��7��#_�O�}qY��[�&p�C���6�Ǜ��X�X��쏞}
�Iפ��{�|F�����:�!��ir7���Ǐeq^we%R
\���h���-^A�6�Э=��n#�N�Ah�]�6'�t�^�R��x�<!fjU�X�H�~'���2��i3e%m®t^^9f���R������SJ��I:R�����=9��RC9Y�Ûl��@Jciy��NK�Πٝ���>Dq�<��|���~x��0M�W�LGz�T��Ɍ����KN�x[EiL#.��Q�u;��PR~�OMR��� L�f�[ƒ n�VL�$FC5�#1:h�y���c"����/��2�Ot�>��!��G���H���Y��J��u�a|���Y)�{���׹=���KĖ��q�FE�Qt��Z�]Y��'.�.I�ؓ��G��N�qJ�zft���4��R��g�	�D�t�PqJO)!3iK�Y#��\CH�H^�F�$'NvX�G�)i<�b
����j4��C����>3Q=�Jt�sd��<�s�E$�.)���y�bV�&h"-�{���f��
1B5�������V��H�tK�����J��Q���]���P�,E�����/6�s;)�WD�K�t8�o��t��
����_+H�߫��ኆ�0E��u�H;1 �W-����g6�M�oZ]��FsF?{�g}�F��Gdz�s�G1j`�$B�(U	�S��Q:A>��na�t]@�X������+a��%�Vu���[����ni��*��QA����-謁�c@%��`:N$�չ��� �G2
�(�k.�
%��/����U�#������Q�Q�ɠ��M)�æ� �Q���� ���&{��֠��y�J�����;���\1yC�q����'d���S�dd�������S4$5��Z~h-�q���`'��+����08{���+�"J/�,*���Vl��*G���UW&sr7a�v
�qѩP���mS�H���0���mܴ��'��hM��\F*rj^��i/����SXΠim�T?<C1Z��A����d
��ؒ��n��[����#/a[_�LCҚ�NaQ٧s	�
rOj��#�"�P�eyAN�mXW
�:w�r�6�{���~)c��-DT]��3�?ӷݍ����+@��$)��}hn���)�c]��A~�K�p��y���|�7�l���.�|��H�=��~�U�z"j�N�&�.h��H�8k�!����M��sL˒���U�
d�ݭ�R�t�C����Y��g����N\���s�"~��'��}�@�F�P{�	�Xs���`O,�Ma�����i�mG�^�� ߾����.z	���A��o��`]U�4�G�1��!����
������2�����!o	,�ڻV�m��g��j��dV�K�'�j!��n�Ɠ�m�D�Ø��a���8�N���c�ح>�a�8m �I��ͼR���<'��}BD�E%�nnB���O]�%No�Np��&#5U��v���~]��L��}���FF���� ��9�i��J���W�.���;g���^���ƬQ|��B"%�HU�HXU{�-U��ϑ�	;�ET!�@���!��.��g�j`�^ӎ=^�Fc�{p���!�mv	/��zY������G�D9�ړ�N�V��,=~s��L���\�����|5"��!��F� �2����?�k%J��7 �C�(��Bh0��zF�#*&Ld�>�3U��k�z�4�����K�rW@Üc�����k�C$�׮�W�\��lI"q ��� E �
v0�9�:�/��C�[s�Z9�J���e���.�F4�ǒ{Ә��,�?�5� ���!��i�̹Ɂ3"�v�\%�ޤV�!��5�g�Y�l��@����/�$����a���0^���u�gm9�"�j���P���b:�O��
�ds��\�z�;<����#��Ы�D������;���`����8��s6.�Hi�k�i�>R�W��H�`���"X���cTk� L�O>�Lb�P&Û�4QOt"�y�C��%m���pVK������=���������G��X�Fۊ}���d�\����i�*��W� �r�X��ř0#ht���N܆kc� �*��Z �a�?���1e�1s?A�z���ۑ�Մ�d��M_$8%2��?��1�-6���2uDs>��*ӵ<�#�&�2>��~�$?ym�i'�g�����jڎn9g�p$*���Y���G�
�	��(�R`/����A�{r��N8�MS��gh!�V�:JY�s��)��������U�:dp���¡9��${ו�o�ywT���';=ɵlT���x�����OJ#��?�j�p�oW�5��,��j5��'Uኈl9:��"߹�(�1��J�>6ڿQ����D�vﾴѴ��-�f�v^�<�F̤�LLA���2`@.v�pm�%ն/zW��ms�h2���]}��~�2�d`���0��auI�Σ�],b=�vw�5��/�8�J�#
u��S��K}�(8m�V2����a��a����,��)sCz� ������i���]N&�t��*�Q��, fXK3�����TA���4JGh���)l*@|�M�{%�0�[�ΕK�|�H��j���D20�!rK��ޯ�*��r�Y=�H�y%"p�tm%���^�<gi�I�!��KǇ���amT?W�Pl2JT �@p�G֝ph�}���{�>v���K!Þ��[���*g���/\�CSUB� zںK����� 7��9��6�(���=R�I�Gk��6�V��#Qa��t�i��ɲ	a%��ndt�ǔ�u4停�Խ��_y��/�p!5RQ��;�YS�~������f��˚ٽ8
�VA::
�W��T�\�`ᝯ����3�a���׆�!K/���ф)#G�%O�))�ݜ�8J`?�� [L
m�A������l�Q%
t��hsǏ�-�on�a��g�ɶ%��D4�~���<O����	.(D�w��g����~�� Z�aײ�A4�+�c $h��n�����r���l�R!�P��ӄј)KDr�������G��<J��-q�HH,+vbAW,�[dzk܇{�x���'�ր�dYȬ�*���+�g��t��ײ�2X�n�f�7� iQ�E)�����.�VH��DL�QNR��:����z�v�C�2,��9���XD�>b�|O??�=&&��~���?P�;��qc�z�Of��(�f,
,�9�La����XI+G���ڭ���,�������XsA!p�Ӡ2{70��??u�ù��v�K���W���VL�w�V�؆KD���΄�8�������¬�HpƮ-�ub�V�����__�A�./��\t+�`�Ɔ )��2���[\ *3(��հ�����E�ny9�@�h��'�;L�h�Y�
�w.(�X3�|�R��O��B�ۋK9�`5��!�I�����*��R�si��r���c)3hOi�N5I�'v(���Q#�@bk������T�(Ԡ7��yx�TP�?�5(�)�0A�n0�8�?|�F}&�,�qP��m��Y! �^��i$�[D~V}�Ȉ7\vz�-�fy^��f!���^�7LBl��yY�\�i@�������;�6^��mhl���8o��	�7�̦�"��SFQ�Ey�����?;%��D�����i�Q�${.f��h��=�o\�{�����i��8;����.<V�W"��&JH�lʝZ�g㣢�qy�B�P&�~�����h݈��@�n*kX����WGi�숋fystp3OVP�/_3	;�nt��l6{���y�"ё��Oة8�D/ʇ���2T�a���>XA��,9n}���C���ж&�4�����Y��Q����ot �ou[�	�S3hKa�v���V�*3���A��Ѹח�I�l 	i���8��)-4�Zz	8����S�'@X�.GQ⳴�I_]�Qb!�=���;8 H- �m��yEoYO�6g�� Ԝjjo&�%��ǔ����
��o�&͔�]�A�M v�0�P(�=���u�L�򅊶�������&�
T�"E��e�-WH?9D3D�UW	q��B�{��c�~�4��:��)Y��+ٽ�qr�3M�� ^X�E��6��`���O�#��y�>D��sC��}z'���:X'�pI�ȓxUa�Kۻ��9{i�'���_�ZPA�G9{X��Aӓ`C��e{N=���0�G��|��L$q��l��ē���{r̐I��!Ŝ���߯�h��x�c��.��3	���j0��"!L���
��t�5��߲A):�r���X��\�bE�uP9�՚=@��}nK���SЊ�,Q��3G�V�e�~#��Ⱦ���h��]9sq�@��[���;�78�]x�*x�rS��d*{(j�5��<T�Ե��H�	V��"Z���f�ޒvx�Nȟ&������Ocy��'��7b�Z�gu*��o�qCy���Mo�'��b�ab�V���3����j�і�DQ�ƽ�܊�/H�6���<�c�U��y7�=���9�������1\<�_E��jnH�O��F����߮�d��uyDe�M>MJ͋����3��\pn_"���[,{��S�SO��,d�Z�ҟO�)POR�l�4��!%�/h��;.#/"Y;�]��vt���&�#h �ǁ�A��I������(	m��؊ҤGޢ3�E��/���?u�+裰j���!�\9�&z���4����~�6(+5!I�, �)�莉C��A��ƀ-���/>w#[i̍6k^���e� AZ2�V
#�"�����C>�!��+vu��C�2�[��d��ekg��'�}��?���g�V	�O������2M��`柔�ע7��+�d����$��U�d~Z����r�E�ex�~I���y��$̙�m��?K�b=�h����uR��Ms ؎k5�^s_A;_��:���B�GCW64Ⱦ�I�uG�c�yԏR.��8�r|3u�u��}H&ti�1ņN��EA芙^�>a�o
%C�еƪ�t��f�[s�0?���h';��!�v�~��!�{��&�`ԕh˥W{�8*�k�T�!5�}�ӆm[vb2��B^:���ɐ*c&֬�B��z���,�B����]HR���k�){B�Ǡ6�e���>*�@����B3����>�x���UF���|�0s��