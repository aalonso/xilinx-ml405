XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����q�+�S���1���25u.%�yk��c���>�*�>Z��.��GW��ɯ\3s������X*��1�;��Zu8 2��:��V���5�
=3&G���T7.0in ��3���3���2' чY�A�z��Y��eb�E��糫ZɓE�&��qi�n�����sy� �΂�{�~���O��^�wd�H�3�$u�sx�F�,�a?)������;ʨ������*�[��"Г�-Ca�FvD?4.Bm߶��t��_�_�[�/�V\��e��"�A�Y�R�5g(����Zy��}��MC%��ɟ��,w����8[����	8P�8���k;Ǯ�P@v\��Ɋ�fW� �X�v3�?'�h){0;bh�d���ƽ�?^=�if��!Ki�2r�KEtywg���KI���1���M�D-�vʇ��݉Ϡc#��:N*q=��!���y���
r�G�ݕ[<�V�2(�V��^͠ y:r����6��%7m�)�V<kg]�D��+W���Q���M����	s΢:�?L�T+C�����u���y���t7�z�:��"���#�f�Q�fۊo�y��h_�:����.Tg��B�r�c��Q'�+�N�9��]Z�Ha���[y�(�V��:���ֲ�Tr�X{+���_}Ąo2��5⻓Y��gں�C���1k����iS
��=�-ַ�¡�a�q:q��;��������N$�.5ԓf�W�F�O ��'ִԠ�0XlxVHYEB    1017     680�Y�QK�&4v��o��/��/f�Υ�����G�v���κ�(厸��yH<	a9�Ǿ��2�#w�}(F����;%Y�����(�H%Gd�sM��w�  �G�����w�M�~6+��&�{�O��Y�^��=P�V��r�n��&�5��f���ٹ[���NڣF}�g��bŗ�� ޕ��gnOm���%�C�b��%�9�.W-�Q��M�eUi�����X�w�B��Ʈ��^�:�����7�Z`p��8b�����w�QKk��%"Ϗ���G ŤI�?��Rv�w��O��6h<�3+��L�f���:�����w
+RQ���iH��ծ��OH�ލ�e����1�vPʏ�{t}���\k��A�B�W����4[��~\I��۪E�z��RHR��*$�����yۦ�k�`��F�+e9~\%�n��Y�T�`/��A]*}��"�s��Ni�0L{+*-�\*�M�π�L��O���)����E�٣3� �=a1���|/� :~Z͓[��jg�l0��]&d�D�mo�UQ��%DF5�7�T�>.�^r%�\Zv�����EK���+��Np��e��GEIv���~y<����H��?I���Q3 /��[���o�CG̜�f�.tM�m����M���2��\"d�aX��XT�°5k��͂le8���~C��]B�D�����W�"�/���l�(�y�q�27���{N�,k�E�9���iݧ���Oջj�>�e�.���ē0�}�u��W�~�.��/��-f$C�P�!y��-���ƚ�⿒C���!r�V�)VsY��6��`i�C$����cIWq�����(���o���q�I�+7�`4Y_O����"gJ���^@8[�5z��K%�d`j��{�$�'ZV}�XI�녃���ޤ���%#t�����qg��@o9Mo�b������?�M�$ه8�cԣ-�M
���p\�B�ۺ��IB����u�ӡ&��+V�2��� ����}��v$�����s�%0kV�H�P_�R6�[�v��+�u�ޯ�2�_�N�N�! ����@@x�S9eJ�����w�s}{B͹,H�}���� &��I����z�$���O�ܚC�ҫ}�6|�'"��(���y���wJ��+JSJ�ߧ\�(�t�	�ܶC��,���%��C��#����tF:��@-	P����5��
@��� or�n5cAx����ի-�g�<0���Z��U��Y���J逯g���	D��r[�8D>�I�E������]ԯ�J�*r?�U�1Xr6�����oHu��R|ָ��9f����1
ON�NG�LI��q<�/T����C�xqrn�&o�b�2]���M.��G�?�oP�X'Ӯ~�,O,����܉�4�y0g�;�俿P�!�Rig�&��1E}jl?,I�z�#�v�߷�,G�I�؋��P���ExY�o����)ۏ�-�S̆0fM��+�yM�ќ~!J��!��'���n��
��3B,����v�u_w�Xi��:L��R(W�@��>���{t{����~(�{�{c\��?db|b���k��_~�r>�cҭR~OJ\a�\�}H3�6 3��ǁZ�+I�b