XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$����U��i<Q+��mz7�@�p�h��&�% S�q!,��V���J<�:縬�����ɮ���h�c'�w6���}��oyZ]Ӵ��
?��x�<�1J�etV���9�s&�V2�z�P�o�0L�VF�WeSC���
&c�������g1�Z3����sns+�Tt<'{y�b�W�����G�f�����:0��N�3Z8�8Cs�M
��M���P���d�6�u�|Y�d|[q�R�T�5��z��i�a\��;��E%!q"��I�@�CxH�`:.k�vA\4�{(�	����*�d���5��)�G/����gZNl���Ǒ�����yH���6�_ͥ�PJV�U[eiP��:�>��:���^Q_+Y���.X䢀�ui��ɛ.�q�N�Z���Y�ʸ�#=�����N��|+��t��1j9��%݆ԭ �#,,@�<�3��1m�tф$:G|���lQ��E�%"Q��U˘%�@�/�$ȫ��=��׬��Kǰ�o��0�XK����3��tl��
��E;#��~lku��#£hoxZ-��{?9����>0T� Wc��nQ����2H��sV�Drz7������j>���'�eA�nck��~[C�X��߈F��Z�w~C�����mý����~�F�]ਛ݃@��uy'h�R�"�D&����	��� z6��fg����*fT�����,*M�Kzo��W��-�1�SZ�3�zrG�L�%?�@%��fgK�:���"�����XlxVHYEB    3e0e    1150�zEa+`t�ك#�1~?��p��2�J����u˴T�x��E0����Iۤ �X�d,��6�>)wP�T�7�2~kv�,�t� Y ��F�B6}ԍ}9U�WQ[56C�}��1� k����ThSZ�`�*!y�YS{b��Bx��������H����d����Mj���E魎8ƕ��Y7�
8j��ۺ���w�x~��~e��+��!*�&apG��W�ba�p᧨گ��橓��R9���>oXk� ��w�@�N�EX���
����8ͼ�#�5�����a�[hY`VBj{��f�\���q�r���J�݊8���P���f���O�u����~��hf,�_�tR��x])��as=���/����O��}��W��-a���?4AP�'�a\�r��`HM��S�/�����/�w�[�)_\�h���V�'�"�ƈK!�h�I�8֥���1�_61=�޵lh6:!�ȼ7P�-dZWY�܋��׭`ы�����v�}���V�0 -X��߇
��s��Qܐ$
rȩP�#���ϐ�C�Fz%8�$�'�Y]��ϲ������
��J��o�:/$�n�'�ட���x?w�ʮi�W�a3��tH�R"�����\.�I[�a�1VX���b�%��y<���%<V�����YFYJ�I�1��_m@�sb&��PLS�*Ʌ"#��j+�ݩ���m#P����Ҵ���w� �g�}�A���K�|���t ѹ|���v&��HT;^��V	4҆�K�#ic��HM~�wL�0F������:�&�X�&�@v"2�
%;���-�{M��7����%X�,����t$O2����$�1�Z<�7ٹ���FZh�C�K+��]+���ݡ�aE?w���wI#�������dMư��@�C5ّ������kg���d�nM��*9�X���W�y�{0b�~B}���kI���:�釰^�p���4(%R�M�ƣ�����e��Dd���V��b�;�U}D�:_��vU�C�	�e	�3�AHY�v��x�ݣKB��*ڑw�Aa�#1�
3���k���puy8����3�T��H�dE�L(Ǡ	�I�Xu�Ea��4"1��CGsD*`Aʔ:�����K,����O�_n�$�J���f�}��fN~!�c{P�g.&�D��:0�J`~�	�Z$�����H�4M1q�)�D#ֵ��sv��%���&93髰<]=1Ԙ�e�G,D���.L���I�<_z���Lo�X�Ӿ��1=8U#�@f�c�[�"��`ˍٲKh$�de�1G˕��*��l���}��^��G[�MѸ�G��AD��Mz��[��&iw|�mN*���s:r�f-ordg���3�������ŝ�N�:m�U�A�b��������8!V�~�8��D�!���J)���{��t��(���Ȣ��Ũ$�Ĳ��u
P��P����u�M40W���{��5�y��ه:�Ӥ����GޕB o�U��6;~���r�G��G�ѡ�5�J�V�[%��KӴ�AS�F]D�)��Og�Z<~�� ^��ѻ�M��0a).LZ�oJa���Hӧ,�`Jh���>�kb�{A�1;��]i�/�G������n̻�u�P�~�ݙ�ʺ�W_Z�Mj�/�F�/;l��t�J�8�.�7�	}k��1#矝:DAE�Vd*陏�c��jm��B}ĴKgO��փ���&
X���Q�'��ȥ��8�E,�N�f���h-i��ga��|7>��6�ŽH�T�<���k������a��ȶ'�������:�8r����'����G�ȽOY�|ս�0��5�(٦7�z�����o���/��j��Hq���3|lB�1/1�z��8�2����Y1K]&]�~Cw�`L����/��:L�~ۗNɆ&��v�5IV���N^�K8�QsG]OrҏuJ����o0x1+�|TL����sv��_�Jl�G���Yцƃ^f�b@�{�X�ĺ�u�I���ԄB�A��J��a��vU�Kp���(���(P�h���)�tT�K�G^tF_�*'������;�=m,:�}O�@Ö�0N/�y���J��K��=�)�2�c󇰪u�6(��a86�{������G����q��CW��j��J �D�k����h�y��ӯ>���lZX�s�B�*C�4����bUy��~B�T����?���o��أ�Ya�k�[��M"�4��'���ZV�j����E��W����/�؀���[�-�읖��`/5h��R�]��3�6]���������uy�!J|��?�@F]�L�m�C�1o��Z-�Q�IW��q�t�����+9M���F#q��:��v�-��{TY��-̭oZtl��ۊ�Ul% �pJe���"�E \O�P�9f }����z�b3�E�������ؙ�|�ԯ�npF�V���&֩y�v��@���A��F vap�
�;	1(b�t�!�S���E%��Gdve!z�Cm���4�-��=S*\" ��&}l��Le�-~�4g�Й�GW���l���?�C������V��u�!�oO���O��rݴ�6��C���OtVk��Ua��Z\3i�i�k��a�g7�ˊOq;A�hO>^.�4TA��u6�����@@�,Ǳk�@�c��|"i3_ʙ{�?Z�輹�`+�y�;%NE�}�7D����Ų��U �)���6��I`��F�DZ�Wce���FO]�d��D�rF�e}�����%Q��@I����b�L?�>���E/�L��K�d���4u�9�-.N ��B@95,��z��=5����������e�ġj�/6�\|&�x�uN+VEC{!�E��T�LA���R;p�#'�mF՚��S!�',�?�0��+�8���B�����\}�Y�Q�@���U��?��UR��!�qL<j�[�V(�?m�NGg�?i&S&�|v[5����7�=���� NIW�E���%V,�ia���𾼮�j�8=f�5�<_�<�%�tB�E�ú9OJ�Cõw�_4<�A,��uG9-���Jt�>r�vl�Ơ�ܗ����gw詼��l��{�=��q����� �nF�*�������U�$�3u�F��<{Ц�ʲѳ�ƋJ�
!�²��nr�L�����!Y�-�e�pK�I�ͥ���j����^�O%
��G��l����k��N}���n��&�����zR��Jp�@Q��~�����z.�z�Ф����N	�3%�*������N���Vv��M��^���$Ls�>��~�H�&t ��!@����qCk_�*���-ÚtX"��a����K�m<O��a��@H��y;����µ���,���I�kCS�"��v����'sa�+C�4�cιߢ�ʤ��ѝ������<��ÿ���	3ۺ� fa}���pGI�rY��0w�/���U,�1^��}��5?��N����G�	�S3p��|^|��̧^S4�}�2	/�B^$�K���AKW�i1�%���i��a,�:a�6��X9�$�+���a���A�q�=���š)��o�A~s���cl�)sf!/OP���y� �"k.�L�(�?����C��+�k[�� �4]4mب\ˡd}>!åb ��eND����wK��;��-�5�a�O*�#0`�ˠ�F����+:7Jp�d�J�J��,���2�z(���KU^����\QR2A	Ŭ�0(�s
�`>�({�T$G͉��WL�x\P��蔦6;��;&2ĩr�ضEh�M%\�� [(� �%Lh"p�_�(^�iLCr�,�F�����);��j�#�)1��.�`C���3>\�c���UTt�����dF3B�l�S�I]����F����!�f����G��dZ�O-��AЌ��01$��J5�z��[:��i�@��7^`���j�.�| �ì%��NM���>�a�6��ű�jz��N�:ԥ��W��V
��8�D�w���6�׼��'�%r�A�P>ր�E( �N*弍Z���̊]��
\�P�9��._��&��	Ҍ�d��W�̹��Q+If��F_K+t6|�b�G�u8�|��s�ж,����9�r��pHI�����z\�iD2~)���xמ�?��}��(N("!8{lÁJarS�4sϯ<�/��"H����$M�U��f��#s
��Z��T�O���n����;.������/�� u���B�`�\�vViɈKiK�)B�����N�,+�h��b �L�aZ��/��H��}����!���Q��Qʐþ��5��i