XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v�n��`�n�!	u/|��ϸ�oꩴ�>���Y�F	֠��2b�P���n���z�7�	{XL�k�+[hE�T����}}�j�-�)���J@��J["�H�úC%��A��t�����NV��϶9<�|^6	 ��즾��_h�s �g�}d�~x)�Y���Qa�44�frM�a�|1����U-�Qj�ZZ+㠦+�f$�P���<�/o��]���P۳���{�5��-9�k�݄�*�š���+�?���ɹ�>}ܻ�J�M�F<�nN)�!��j���#t$�'v'\0�h��Ǚr���	#rYC���$�'�����T{EY(3{�`���x�X��Rř���L��{�V�~�������7���
\tN�&keg}�nJ�����LW���L;�ɒ�� 9����<y[$�i��}1����F���$z��s;EsI!dȇm�����S�u$��<T���[	R\vY�Z6���/�HN������:o����L�~y�C�*�i��2)7̋��z� �h։o�O|�hr����H���:˅����Z6�~L�£+��8�W������I$Λ�Ղ���5|V:��E�q�ݥ�WAlæ���=ΰd�}ϪƊ<��g"�Y7R�$:Y�V�ӟ�boi�iD�v�h7�!4lG}eҠ��q�Q�>�hƌO�6���L�v��m��9���T�{)���jޘd�����ƚf���$�� ��?�����������^�K�^��b0Ճ`�J��I��bW�XlxVHYEB    bc57    27e0胪�:V�9�>~G1��16��_(o�My�E�z)�,��0
$��,z�LݱW�ч<�6�f
m;�D@�x�d�B�xI�O�0͖�ώ*��O;HB���S��A��92)��L,�JF�X����V�e��O��5�p�Zn��T}����'���կ�8����E���nhP���Ü�}?���a�yX���M�t�sl��	��v�	\����7�/���ݖ�\��J��l��Q���#;Zs)��^1��P"�HE����)�� ���ڦ�o�L_��.)��xѕ���~���_U�G=�l��,l��4i�����-�^g��Y4�������}H`,Kv�*/�Y���0���F	�WC�Ё����z�\}�8ʱ2v��=U���Dl�M�7��7�{��Vy�uXR�8�b <i!"ݰ��C��Qf��*��vX|i=�2u���&��ܛ�_;��z���[���UG�lyQ��iӀQb�b`����ۙu�gd�D���S�����=�3$��x+y��eK�]�r���Is���Ӳ��ef�ϐߧ����T��eA���b��:J���-�<��}��R""5't�0����7�_IN,x@���V[�jIs��� C�I��A������&-�ٞ+��N>��@]b�+Ĕ����k�ŉ�Z��<X�+�P��M�{��{�]�ʈ��p*�R��b45M��|Ծy�H|#F�.@S,R��fY�}M)pi����<j�3�Mx״��%���_y��Z�cBR����]�-4�v�2����\�J�͆G�E��uY=L+3^2'x3�!w�r^k�.��{��h���$r��aX�J��&�h�����#چ�EG�o�#�J�>�%��{��QJ���a�����+�ʘ�L��R����&S���.˰��fR�=� ��i�A�O�jx.��$+u���t�_��N��݂�3E�Z���TS���+� �`��UPOAt���fCl���Xm��y�PC�w-.AW6�''7ǵ�Cn���ps$�0
�3<��<[7��2]�����Kk%��0���М����0x�ߊ`���#���I��n�<��k��O������zvϺ'�+��+V���	��v��1E��[r_�GE|�"g��I75�AV����k�����et�
�u㚱�y�6~�B�PEp��lƝLH��M��2��Fj���#�CƾK��׾�s����o}��%���ݱ��+5,�#aQ���-j{|�a^���)�?�li�hֵ��<��Ϳ����C��3{6�����̈�/����&�w�r;'i�[b�Fޟ���>_�fHu�_T�́`�@��O�������+=	��l:��~�0�����g���7
��uJN}qng���?YԒ^w������E���2�6I)]f�]ߧY��7,]�~)J�,`}�kb}���޺�<>p5�-.ឝ�TG�;h[ 9���xrn���q��.:�x����5�>D�h6[s����	�Q7\�b��;d����m�ԨS`ө����(�#0��B�ǁw3P���R��n�馟y���_$�?��e 
[�Fu#Fh��"�8p�0��ễཷ+I&{]*��U�좵��hm�"u��7Ş��8=�6�)�49�T��4~c��	���E��s@�ھ��k2���P�d-��"���Ƽ�%����4�8*m���
��Q�X�̝�����7X*�z)��}񒣡$����0^�E�i��̶��j�p��y�_Yy0KN>���
�/^*��r��8Dd��6�܆�6���:V����!�����71@�|~�֡ijdݓׄQ>��-'���ڵ8Y8ܷ	.R�4�����Bt������y�z~E��8�u�N �c�7�=�*hr7L)NuԺ�|���֟~:��~띡w��t�����k,l�=�"|���e艱򘖰��>*Ƨߜ֏�~��K=�ͯ�(z� IY��_�cN�0��vLd�L��$,��|���E{٪��9���c�M��g�d�J`�T\EC��i\G�,���jh�/H�V��O6,�T~�Ik_}�ߟG��� t�P�I���bSu��\z�ŦC]��廩�~�޳���"k���$1�_`uP9�l(�ӱ`�7��d��]�"����׏�J[�߮M8�O[?*��}
�ꀘ�O�DB@X�%�M��h��� 7z�J������!)?~�̳nk�z�h�&(Y��7_�����9FŅ�{�3��4���Js�S�0�q0kOY(x4v�t��x�h����/�����V[�C&;�P61B?o:n�T��*���"d<�r��v�C|��G�ʄ������w������)����P[)p�)T�i%Q��ʣ�]/l����\�pUi������f��v4��=d/��<k�ىLS_���$�	�?d�qM��mb?Xr�1��g���'䞵TF�Chx�a��f�-�4�����KUɰ�U�tmW��J f?ҧ�V��?���@5�b��!ƕZz�,�׎����#z�Qژ-M���7`���BTꛨ7/�դ��|[��6�Jm��,�c��:�7yh9��Sz�^��3^���<�����*��I�$�Fq�Q^�i���S�.0�B�vZF��}�,��o�)�J�a��J=\���L����e�Ϳ"�K�����;n�)*���m����=*�t��,�O��������E6��/eK�����ʗq��)��bF՜�8Ev�[M�h0� �?㤱��R]�
�Imd=]��5ɮ�Fz$<��yXo~��<9�{�]���� &���q���"�}Xrq�B2P�:q����/��=>��M$�B��eaB��<�oA�S�LJm^jnӆL7��n����C+V� �${̭�O_�/�vTT��$v�O��}1V=�l��o)�WJ�;5U�(�_�Q�ӳ����b���c�4'�Dz��H��΄��#����b�sOPFn�:���i��	�O���'ٽk�.���Y.���8}'���׭�e#�T���� rtx�b|����1E��1�=&��:@R���	T+P������[Ds�����"���V�����oX3�|�ӯ���ҸUI_�Q�ϫ#��=��L���m�
!���a�%_)��:������?[��[ٮ��1b�.ј���5�8X��}���Q~���\xn���+�Ӽ�*��^çX���v�ާM1�s��?
�e�s4�։��J-��+���J@'���3s�K��hAzͣ,�ӌ#�'#�&�j��#e�;9��+�ݳ%������kk3���5�'N�s��+��=J�Ă����F!z��җ� Ieb��G�lb�=��X��4/��K���K�y���a� �R{[t�[�}� �z��_�1�B�xcS��{+�9�}Gn�dً�ϫdRb�39�l\1;�&7��+tC��[�k���� M����	��I�1C
t�p5�xZm�c~�c�ؙ����	�Z|�<��<���q��q��	����gӡD���vh�A�N�[�8ǑZ��y?p��Pa���͟�K�A��~�D>�}���3�A��Xtn(�1�Wɖ��Pk<	D�(3�����|,��^f��Ʀyv��wKkT3v���죄���3�L�����/�b(b����zD��[�-I=� ��P���x#��Yx��%`�:�G����F;AU�$���ص4Í�!('�l�4�+��{��:r�Hz�w�/#4���C��7|�X_����R�c�U�^���9�O�������H��R��۰�̣"�gB���.�&��h䑖�D���RF"��/�Dg,���m��'v�� ]���#Yty�R�m3�Ǵfz��V�	���O{�O��i[�i1�u)|_m�K�c��Y�Qc-�F�8=E��W���&!���^N'��蜪^�k�1�.�,b��r�)�
x��$m�����{�߳�%h�&�%8ep��������|���p�AU�.�Cq�����㠚�y��pV����^Su/)��qk�X�h�w���_�a�o-�Q����Es�H���ط��h�����whn���Z�u��p�}�' 3b��5��5���}W죪�Z4�gZ�ب���?�SBQ;�E���_� ����h�B��$�����Q�,���	Kw���rn���"�����6+��{�Xa�!0f���_��x7i�;������_lxx�ƛQ-�z�^J�,�.GQ�Ý6U��b-;`u^�e`>]W::�7�Ԫ�F'�p�*и��
/R!��o�PXu�q�g6�g*����1\�h1�_.�yQx�q�ʅ��V�5�O���0��;���N����
��/��ҧ���F��.����0�`=�RiMA��c��n]9徹;�T�}�>#ӿ�7����G�%?`bo�<j^�Ҳzˎ��"cMN�Azz!m���zJ����L�c��� !���<#��I-�g�z�ȗ"�&��0�Љ�����&`�x_M�]Rz'E/�!LF�~j��H��y���h�{<�΄�p�vI����Ȏ +�X{���V�=�B���W���B��'�2�[�>.ב�)$j���Z'���ۖ]1ԟ8���Zܱ��	@Yi�g�`%����X;G:ܗ�Uɯ�'F����I13Bv�jԁ�k�]��& �%ny �
%��|��q	���G��������54�+G�#3s�{�ާG0sEU�d�k?1�,���|ج��'��h�m'��%��O��=�`�ܶ�dh��W��Ð���ϝY��!��t��:8J'�1:"1��@v�lrW�F/�N=�Q��@ �?��K�a�e(�O�G9!�57����_�qx��0?�gX�7�X�@)7T�"�@=���g�)�5�J���G��
�9���P/�����i�W�4�G^������Zr=,�xl��fIۅ�K8����]������I���)�o��q|�L�rqq�Hw�m���n���֬�]~��l:��K	=��i(F'�z�]z���Q�����w�.&�j��Й��D�Z���;���f��zo�t[<�o3�������d��"⡩���]<`m$5����I��!�af:�g��WZ[��8�Y�&�X_�,�P��2�K�Wj�>B�S��)�ǌ�(�*��b;�"�����B&IE�I(����$�^�������b��4��<WxLf��L@0���CDJS��� ���9Z� ���	����xzbχ.�?`)�W���w9��9�e�D^84���w��i����%
f۠e�m�	�K�捴���T�\�9X\p&�yU+�X�
��H}惾�s��H#=�H#.?�{6��c���:����}Zu����.� �ϮQ�䧢��*Qm��z�i�l���'�Xf��P��b\�0?�ȭ��ݩ[�h� ̓6ì��[��K���q��Gտ��r����>
�3�o�F4��d�]SEa�;~�$#��VJ
t`��ЗX�����UvS�9�+�-) �;���t��ů\�V丷6�2x��e�]?;�� �5>K�BM����3�	��=Q7���[KL�)o1Ï�����f5G©0���#�<~h�j;��)͙�_��ti�zD�5����	��h��ҹ�O2��S�.�x��e�qk����E�w�(եн{�UgGb��5��ɷ�U�W�6ͭdR��[k�q`� ����=';>v@?�_q|�t~�Ce��8G>fH�%�eY��Py�:�<�v��@P9�I"��s��	zn�r���=Y�ё;�<6���L���p��c��u��Ro���ҌE�w!V��G��s��yJ�h��U�u��T#4	rQ�5*�H|u�(�:���ޣ=� ���-�@�.�c�@����a�B�b�dO�x$�o-���ɢv��齣@@��c���e�ڧ����%�o�6P�!���0��^�w\a�ki��1G�PFr�4l8i�4-t�R�F�9��h���o��Ln3���'�f?�����TA���?��?Z��+��3Ҁ����b��l�1?�>�g�G���^�@&%����T�e������zVTp�~����߮�i%k}&Y�4PK�>���g�l�dܹ+�@ �'�pA(���{�zи����r�19?q���D�˲���&��PCc��@�x�� �#�xs��5�E�q���c�f���Xp(h���zA��|	�\)�=U쌣�����3vVs��j���o��ғ���V��P!��IU��8��!6�o��̝����x���?��[�B/�B�u�T�J� �1��h���S��Z>�M��uoU-�<�rN���/�S]P^M���C�)��BAD�߁D_T���E�����B���ѱ�O��͢�&�;E�;	�7��/��_��v�������.+ߟA?�AF�m�i�m� p=`�-�y��G�5t&�2�4���H�sis��#⏽�F�5��E��k�֢%����-�L4�U�n��Tz�N��p�J@��,R`s�;�xݼv�U�~��v���e�%s���4ɛ�ܒo��
~9� ��T���шf@=
%|i��v3e�xˀQp�isO�
+�#��d����NŎ �����FC���[���~��z<Wo
�}���>�&���=铕k� ��Ѕ\��r���i-f�i���x&@=iƓ5�;�2���o�s���Ӿ�$1w ���&�q^Hn����dy�az�aK����`�Y%���z ����ޝvf��#x_�Wh�O6�\u��\����O�Pn��� �!�CƓv�G�:����t'��`�9��]0U��1k*!�i�AW_�R���k��#k��sP%�Lf2�2;%�~~q�º��e���O��@�u�	�(͠�[�v�JWo1�1�3R�n��;�N�nV���C+��3?��EG2q�����"�
��+�a��ɡ\�I97���gjS�\|�5b'�P�gC��|a�j��,�#&�{�GC��?3���&/�x�Fhx�P7M�����kq!tpXn�4[�*�I:8�<	A �A�:���=����9�!|� �wQ��:���o'C� >~�fnM��[!`��!�2J4�ZZT���-.���1Jo
u�K��yEӲb�.��E�D�7F�"�)8ӝ](����P/4���bE��ԧ����m�{�j��F���4nrrW�؂�uQ���JJ���hOF��(okb���˜��-���DN/�'���<�� ���WO�Y}�pm8H�\�ֵ�2~�v����V"6���a����M�����`��6��$��I3�ܽ<�L�7����ҵU�U>�����'��Ͼ�,.X�U���ϫ���D�$�5i�B�~�pe���һ�"���y_�C��jl��'�/�\]*�{OO�6�c!l�mu9t&�yL�����7u@��|�-1eɩ���,)3e�7�ծ�q�.�8�2�^ޅ�ҸyN	���9*[W��U�	'��d�X�+,&��饆ܯ܋�	߬1�1{��X!n7�q��n[���$�NY��F�V*{�B=�$7�������Ť|�"����Ja�)����uLW��W�f�/��>��sf/��������6%q�p�<�[uYɾ�fp�<��Mr��ô�_�!��CO��};	�b���\�St9i��l����׌3��\����嶱���R���R��m\P����S/Fv�¬�}��֣����r6y��K;�:��t"ԂY�,�Q�|;�B���#��2��.g��G�����y5�4��*v��]����㬅�����T)�s��ikJ>+>X�Z�K�2�����[��Xl�R��+-��!\��@��^>�O��A��`�c?�|��6��z�N�z�1��qmMgO�ͣˉ!ʛ���,}�%���]>��J� P0��巉V���,���Q�0�FP�1�W�����<7�J' ����iGj'F6Irz&�'��*9�D6�D����$Lҏa�p��'om++5�k������^�iyn ΋Fd(#pɊ�
|��O��KV���=��AGC.���@����<�J��x;�����9qP�VY�E��S���>V��:�O���bK�cd�&�bغ��#-`?n�y<w{m����o�Rݤ����twm�r�#�Łޒm��l�,���&��qX�<q@�� �������K�;�Վ��ȩ�?O��������Uk�O+8;V3�l�0􅟙�|}i��"Z~�b�!�ҥD��x��UxD����a�3vrd L��8`؃�q>I\�9�"�s�E�<y��o��z9i|@���w���7�"��kd��	R�|���(�*���t�H���B?=�U��Օ�o��ᯥ�w-���T��\^1^9�׆��g ����%@|�~C�UE$a�.�A<}qC!��͜�a^P�OYw��x4��_������m3vW��P	����Zm�(.}7��1gD�*JMt��L�k[^�݆����*�ß�9�}!���?��d�3+J1��� �*�q�3��c�;Kx����@��e����/4E���]�m�P�>Ky�Vd�D��KpQi���y�Cⵁy�6*䳲A �n�����I�g��Q�V޼��гΨ�I��Ecah��
�A$o�)�,H��;YM��dR{/3]m����Ul��G��A:WJ�6g��H4�:�[���U(Lt{�WK���)]�l�R���5�rd��^h�&�C,�$􇐬�Dw�oؔ�5���4;�R��T_涋dI�	zd�c���%�`F���|çŜU�d2Sy����']��L�����Vz+"�b�z{JS��
�Q���]��_�S)966,BTrT@J�9��_��h�>\�?'��^ujz��]!8��T�5/��z =���}T���W�P"�-o�ȴ���YG��8�
F�ʗ����o�\�"��ʪ ���E�� @���'XA�� 93��+9�!�]g�:ي�rtMO��~�ѳ��aCG�O���r(I!|mm]�ͼL�m� �!5��!��e�K�s1/��Y7�:
�A+�j�8�u��c���)8EZ�sƶ�FL��).te�	��?#���ę��3����ұ񹻣���'�e�H�UG�k)�=�	ID�������dh���V@�b�����k-����{�OQ�m߼,�+�q#�����YbD.���`Z
��$��{��SQ�ɏ�`H��\Eg��k��4i0��2$.W&������EIl�5�6����
.F���Z.��}�1�-�����ɇ�J��X�+kbB9���C% �M<��!�0-�/��=��5O	ۈ��6��k��
��O�QנnogE�.Kkm��v�+. j�!S�B���Ř�u"�ގA
��$D#1��ҡQ����ֳ.��8�|'�2���t�xCߝ8���o��O����й�� ���MJ�[#�1x��e��|\1D��.��`	S+����0q9�z���B�k��B{S���&
�w*�f��e��\{�n��Y��
ӛ:��)�G@u}?{:IT!�Pd��+��R����?���m���d/y�!���m
ɺ�Yn�^� ��t��Vm�Qg�F( ��15�/��0���Q!�U�{��1'�E�h�"����߃���X��k��h!a<YA������ݗ���d��#G����Ln�8?l�����:{�;9rD0������Φ�$,��~~֐L�*����n���ȭ��Q��o/hwƚ�:�����t��ҸDՋ>���°F�����]|!�@Y���������O�����(Oq����υ27t�P@���H�Ee;�PX���IP]hä��C	B�e�e�7����IbJ0U��Žs�y�ͮ?�B"�/C!��1a῱�I��M<���	�����K��GM�1�22�x��=L5&