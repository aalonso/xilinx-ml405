XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���*� @#J:��Z�T䅥)�_ШD��4��8��f���E7���Yc����4.�K����	Q:-}{xt� u����k,N�]�!'����ϼ韬Pp-� F�sI�5�K��Ya\�Z���B��E焗!b����t)a]�V��%�����?�Z:�*�)TK@ƣ�����,��w�'�!� +mH��LGCڪ~k�=(�p�/Վ��: �|QE�iA����p���̺Dz�o�l��Ր��QxL��6���7�V��_$l�a����C���Z��T�G�)���V;��*_�@1`1w7���g@z4�-�a�}z��F�4����HLuz�'�������p���������?����R�@��%9��݌��q���u�I�x��b�����Ψ-N^� I������]��&�}���I��?�B`"�R�����b᭡�z _/r�V�Vj���҄���[��̖�/�J���}��O�"��ջ�@؟9�,��ZU�p�	�W&�>UU��5�`2�'���h�X������ߎ�]�>է;&%>�T<=i��`�r�
��j+����/?������f���¶kӎ0�W��6�/���9��9�Xu5���m~�������[N>��#s�L���i׵5��Fl߄��m�+�M��O�| :a��j�4���?ը�Z�k�J�F^�PX��v�]9-���ث�]v����:��zw�!`��ir��j '�XlxVHYEB    47d6    1030}_J򬥔v���Q������L�� ��j*�ař�]�s=e?Pe3w(��H#r-���e�?�%�c�*���ա�18��J���^��}/I+ *r§�f���z4�_���W�G�*��ɮ��W�Z-�fN�l ��rߊ�ٝY�Y���BLg�([�7k���m��Ӥ1��O7u��������10(g�r�lN ��m!dB0v<XO���T���8���mYch�M8��1��Q?/G$�i�X�m���=J�]��f�)�F��[�l�L�N�����ˎ	��whm^�G<����n��a*s	��|������^.��t�p��F4V ����Ӑ �C�X��1RO�:20Z4���슆O�d��OU��I��_#]�9�U�	BWD���d:i��3#4�l���B��)������h�o�(���Ig[���輭ǡ��s3h�g�Y�$N�cq��B
�Q���+��V����<5���֪[u����V��*�נ�5Y_�D��4��^]��P2o�wJ��Ѥ�1@Q'�X��%	�ц��_�gYC�M!�jZ�i�#��R�^��>�wi����+q���M>�i��"��QU;�����-RH���K5L�#����m�`+��1zNK��Cvh������7oD�K["��i��Jÿ����|H\�M����A�uk�*��{� *h[��,z�3(�V;��(K�^�9/�V�O�:�PB2Xw~]`,���M_	m�+`A4H��O��t�\���\..�:��p�jϟ�tW����hV��[iW}<&��Ue~����OL����	�h�]�	�6`�a�o���l���m�K�L>6�R]��&�P�,�m�{_�`ݻ����vT~��?�>4>����v�W���Wl����@ZEU�1���F�v]+#��{�=�ۻa�j���P)2u=���=,f���Z��z���v����wu#��9�ē*���&m��.*������/�e��tbح�������Sx�v���f�6�J1g���� u��Viн����o��\�5�nq��"aBh�\����ZW��?��)�o_� '�8��M^	���(���K�l��%����1/��"��_w�N����c��yi����|��d�w��5?�ḽ�O"P��vx8ot�+=_�
��=�ѣe6��f��>�K�?�a�}���.��UmZkIޞ�ga���.#��p�9e(��(E4`-�]��"#�VT��]Ra1t�R4���+��[����Ɤ�l.ݔ'Xbs<
�s5&4�N�]:��
�����F�y�@�(C﭅5NL8˗��[L9Y��䠴3���X��W���h���o�!��+:_^�'�L��C�kd�b�0d�چ�~(Ä��q^xx�Jsp� ݫ/�]G�5]m���0�7�u�c�'up�2�c"3�hz�ak�<�:0#[`[�����.��Euغ �cw��x�a�`��xƾĆ�_�G������+uF<��n6����	�Ni��	�m2gj�㡹����t�Y�J0�uo�n� `|����B4�)6T���3KTn$���rFM��p�V-�#�PMB��:����"���S{�[�D�F��Ì�Pv���ǒ�N�nC�����ֱ%J'@Z����ʐ�uaF {���C��~@���4���?J�PH�$4P���b�f�����f�e��F�v�U���w��.�R�kwF�u��b�;G��
�ɑ��y>@+��� Rc�{�^|�1�e8���~5j�Kؼ���e�r�+?�4�#���D|�m�,�Y@��0��2���̖��VC��2����	���&r��� 6v�u�O���o�(ݱ])�ɶ��L���|(U�J,�R<u�s�vr���t4��Hۥȱ�Yȃ���P.������<`,��BGlTb���Ue�� k�k'i=2l��3�y��EMd�?��m���b	'R�ɱIH4����lr����9��0@�Y��#UH&�~���v��.���OC���w���܂f�+���-���+��o��5Ӧ�%�[���ƶ~1�9�F_�7R!����}�#�1�g�3� ;�ś��F��7�����IҔBy���Ά�;���Xࠂ�O�.7�y��qL{\���zSAE�8N��ǫנ�߆�,�91	���@�ʌ�'%�o��+�rJ
6HrK��W��ͼ��N��s�8��r\�G��=��޼�gx���s��ٗղ�UPc$�S8��Й�����)�y��O���S��H�H����e�c��=K�%�e�0GY�N�9�@��d_}H�TT����_o��9?´	B�����m�$ȹ$B�$_���[t|��K���=�D���/%
-Z!r�X2��7��媊�m��	w���W�C�'J:͏�j �n�Rw��X�W挙Աh�6O|V�Q\=vc�����Q]3�(���sm�v�6L֧##�2^.J*^�+ٴ?�|����j
����cyY�`�7Bp���e�*W�T���XǙz�'7��]C����!��?c�
��A� P+'ܿ��'�3��j�tZ<}Fʹ�&1�!��}��v-]F�_�0\!2�t��W^䛷��F������0�()�����U$q�.�GmAhC��p�R�L!;���j󋟌�Nfo�tC`��0L����/�y��r��7� #iߜ�w.�b'��8��F���$|dRv!��.BHLxf8��p�,�BC_����g�W��u}�v�Å?��.M�d��:x����1w۫���X�oHm��
�&�
���d0��V"(%�++#
A���CѺ4�(�v�����P�i����>��o���F��4gh2t��5�j q�]��@Ά�(����)�5�G֝�ӻ:{^�����$�5�[���Mcd;��s'4�.�VX��nSf�; `����?�n@ml�/�v�94S`�ޯ�7: 4��4�g��͐���e�Ux���Eb|j4O��n�=,�����)�붭dh`��LD��s�ѧGi9@n��8`t �|2�v��Ӥ-�s6�t�qvr������n,lߝ�
��G�m�ꨲS.�Yy�%��rG��P�t��	Grp$:�<�~@<�}�Rt3ɹdq��|�|�c�5{�������P�x��w5��B��o�,�@�g�CJ�yu�%Y̢G��۬:0	������4�R�_�g,t��ئ���HF� 4l?t�Xƌ�@�S�V�����%��=��O<�g��UH���S���:��z%�fJ[n��ΑZ1n�y�{�S�F�r�P�)�h9��Ռ��z^8����D�z��)�"�8;�@��}���~�9���>�����MR��u���l��F#C���?�^�	�ZJӀ?��U͛
S���G�px������uK}�#�sK��x<$7�떹x��O��`LM��'H1�ɫ��w�o�4~RK�񾧤ݛ�o�ğ��yrx@i�۞�w��b�ˌ`.I��r2�[Q!���J�=��Mt�B"��ۢ<�XG����A>�&��.��!	z�k��#N( =���H*q9X����q��|����S.�I��M���0�)<��u�H�H%��c�t����fC��H�fp&jx]�LpJٽhDR��\�������A6���Rh3�Y�m���=tx.�g,�U��{&+��[L�¯��䕟��Ƞ�[q��׾a���3yM���k�p��4�&����^Ӫ9#�$n�~�7�s�"uL/Z�ʣ2��] @]���;mk���'�%6��h��G!�z��ë�HyU7���U�U�D�~�B�0��4z3�����m-}�U�ӲD�����rU,5(O̠ ����D5!n�c��w^�Bl	U)��� ʭ���"���+��h-�!��-D��-�?��/��T¹�:\��������Y�Y;�!��(WiԎ"7��#�;�� �;�=;��4���'Aͩ�h��ݪ�T��x��
莆�@��ۖ6|Y��>^8i6�G�~��������b9ď1pBh