XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��%S�Ry������+QD[�-y!{��\�k���,EƁF2N�z��b=`k+�g�]�����#�ǌ�nF�S��V����>�����2 e; ��G��Q��D���ws�gkS�濼1��K)��G1*�������,1�]��X�����ARh�V�v���z]E��b����r�90v�qcg$5w����9"�萾�N:E�P�L>yP����N�Uz�h���.ɶ��?�(K��ջ��!��<Xd��oO�$�r���Ϣ�-�Y5k2�]jHO�e���M����8,.=R��}�`P� S5Ѳ�-M� ���٪�j&����j ���[5Y�A�{��T���	+�ʀ��3K��������s�M�H�(+����P����/�QyYulI1��z��R�%�~L�������'{�|����Eڸ��Q��z!�j�=mU�fn��ͬ�kڊ{`U~�F��>�a���~�3KM���}��>M;��:Z8��0'�'�e�N�_uS�tl��Ay��Y�7�Yq�]�V�A��*%z�)���]W[g�بd�?��:G�v��Wd̩����d�]��uFr=���TY�����Y���/��r����to��*X>(�л���-u�Ly���]���k�]KѤ��@���	��4-q.�ךc+��f:���>	J�+xݳ�?��^�S��}Ik���j&�b����[�NeY.A���(��л��z�R�3yd�؅�BzL���!XlxVHYEB    4c95    1190+�-�.C�L!~Q�%�LY���� #D7ŷa�C4��VQf�Ce�%*��m�`;�&$��+?6�fO%��P9o�=�,��|�,�Un[����'��y���@2N�c�����n]rU>�u`36��jh�D��(��2�4ދ�U88l�SfBnBV)��3>��1���b��$"T需���$G����{�W\V����aa3#�Kʱ*#��W#?�l�X�uIF�����#����b�c�._��Sq#��}6Y��ٰM��:u�!����l��(�9��}�:Ua�������1&@�֏���1�-�vX�#�=�ҋs
V>�3��#(��~zxIGׯ�
����0�{LT6�~����]vx����/g5�SV��8&�.1W|zGM�ȵ|�����s#���`�R��[���|I���6g+B7ٷ�۬�����O�N�_�$���r> mAu�2a�8A�&�*`@9H/;�0�%r�iW��?�9�s�^�t�cg��'Ѿ˾�ޥ"�J�,7b��Q�0����OQu�;S!/SaY�ž�z�g� ��ro_n����}�y!�r��zH��_3+��o���i+B��VԱI��g�[_�p\��׶ q�	$����sN��c��I��65���v@��WV��u�=�V�D�Gϡ:�H�6���L�O�8753!���M�GW��W�	�U������M�,p����V��	�x1�s]���9�T��.9�N~M+N�q����
4��V�w�T���y��ߪJ�ߋ�>�����T0���W��b� � j���>����d4)�qG�"�[]J��(\�Ts1���XpKl�v�t�&��z0=7gq\?��Ř6��v���"�	xibY�/�x��a�x�$L���e�\{�?"D��D���'���<��Ci�+-�x;4:���#��Ыï��*�wq�� ���H���F�!�]��[�#��2���=�&i��M��7LE�О%]�w#)<u�Λ�ya��4( G��8��+�/rE�&wP���a }�g�<~�ٕ���c}��ܥA.P�$Lm�F�փ�:GJy�:�7��B�٣�� =�BNFod�xa
_�n�iq�O����so�b*ʟA�6=K��oȲ���	����̃\pO���ci���%Fs�A������q�J�[w|WJ
�3q�>�^b8�*3�y"�t���s��цy����d�KZ0.!�!�φ�!�t��xzc��FV�+8��}�޳ܶ?N oO����evWӧ�:�d���Mw7%1@p] +�}ҹ������Ox��}~bZ�*��g��·�p��/��g&�w
]w��Y)��/�jL���q���N73�WH�(�P_4�EԬ�j:X|M0������\�&� ��ph0g�i�LF��|��+��9��${&�� �q���>�,�)b$y`�#N����R�m�lz����*/f�:�$����ŀ�B9�`�v������S�f�#�H����֠�CQ����}g�iN�k�sW~�nU��XP�5J�:�m��KTb�2�	�9��q,�.BȌ:jLV����gTB�I}�Eԃ{X�>��o�k�h��n�����!���Pd��2a���e��O��f��8�@d�媩*��V����(a���||�S��)W���T��U�U�|+���+Lg������NN�>�Q��YH���cʤp��S����a#����|�'r���9�2�x�����6U�cd�㏹�@^��~[��G�I�����r�^�� �L��1M��f�-��%��N�-��P,��*�b�YO%�b�0G��o�K�ET>@'(T��j���H�:�o����B������GA^��G�������ps}�7
�m���7���fٯ��\�4q��!,��⼪"�IL�s��Ļ�9}(W��%���A��vʛj:Bp�}M�x1͋M3�G=�q��	W�0b�$�|h���H�
黤�K���j�J
y��>���M0�8�`��gM-Ѕ�4�:5V�o�h���+ ��<h�;K쫮�Oi*���X��M�ߥ31n��R�
1O�ٺ�>��IM�>��
��
foJ����M:Ǜu�i�B,�(̜������̀$m��d�8��C=�gF�=X.�_K�����]\�m!*�A��b �i�2�t��V3�t-��r�-i�f�`C�'���HN�^{��J {�2��A�azۺE��=DQjP���r����Fxv�ِ>��Y����_�J��9F��	P�sk�$b��I֖���}
�}ɤ,�AMVQ�Ea#�L����K�v�\s/B�	�w���,�����щ��ߦ;���v�E�J#�o�l�	T�8�����4��S�,f���AU��z��h�E���M�>�3�<�ͧ�<�b��ɶy�J�S7;���MRmX5a��aJ~������R�fD�R1�bX6(����.����I��N��x�؋L�t`+<��I�Ώh9�w� Ѫ��T��-3�d!dT��O�� _��p$$���y��0{]�O9��\��:ӭzg���6������|��vF&��x@�R�t�!^)�Mj���в�5�QӨ��D�L{���1�&���0�9n7qr�����
<�����~wy�3��2#c�Uc}h�AX��K�
R��'���[m�}R��A�"Y�Ѣ�ю���
�a�1<�L�6S\�-�'�2�u���ƈ��A����eE`�>�Y�x��OO�z���$ı�GlVM����ü�8�9���i�x*���Vݪ{1�?4'G��*�8�P8n�M�_��d�'�fO�;����tr8]�E�q��:���	���R�S��1�a->@��emK�Xd@�x���M~־��%�S�Z��ݩ�e��;WwgqX�=ݢ���P�Rw�e�5�x}��,e�ۯXe�C���n��z�y�Y�B	�/q�=���N�uޑ?��SM`3��}��4>m�l}^�!�)'r$�6��c��/Ƥ �>g���?pG���������Y��v=�jp|e�.M@�	|z��ٿ��4���!�Oj����w�^��]���+wP�z�L�0+�Jث���p�������D���,<�{<��ۃ�~Iʄͳ��Q����T��w��qzc��LU��)�8v3�@�T�n�[AII`Lޜx�̦a��蓷�)�_���Ǻ�c��P����G���v5X��%���o2P���O�m�*�o�0T�-��k�䮭0c�=�#=7܍v����,/\���y���1-��� TӞZY}]L����0��c/���PuC=���dx�i@�OD}qq���J��ܧF�47�U��k�!9���>䎮�΢#{JnK"���y��r��6���/���S���촽�t�w�h%^y����y	�- ��Y��!Va�f{�"c7׭g.#��3��)I1,�5�?X�?<�7�@ybIr���c�I��V8���FI���7��^��p�嗿7z��2���K���c��N��n4.��i���˵eXb-C?��#>`�n��S
#8�A>���%�AӍL.M�����:@�݇>k 9�s������ ��
�7��.$�v,%���/��:�d���&o)_PR��
�{	��4ͼt��3���fإ�@bh�/��*)���H��II³%PഹM�j�F"����Mi���"1rs�'��9�z��W�J����1���6.M8��|��GF�B�~�眂�S[�3\�$V�b�����q0\� �[�Bm��ޱ�,y)G�߰7z��<<���;�]�L�g������6�V�O��?�#�A
v��hB7�Uǚi�b4�N��l��%m�5�����#%l`�3%�2��6�g�I�s�"WrP9����f�'��,�#��;�i�m�1G�HfJ~^R�����l�ea��$�A��'"{-1l����dl(l�x������� ���	aɠ�z\�%B��,A��o,�GH4�/���K�=V�����3f�a=�d�p!,F0y����p����Y�4ʪ�e��DꨂT��Ӧ"��S���2�%��`��R
��r.��*��'���G�e�˟�T@ ���#1^��γ�IP���u�{E����%�)l��Vv�
���1�s�u|&������`�4�DU�y6M�i[��� 0�V��%�$��. ����ʹ��1a�.�DYL�������#[Y�lYR$�a�v��+x�Qx�~�{��T'{p5�L(�)�R�i+�5y��3�4��1 �~���w��
~=��7�*QU:��Aۅ>�b��.���V@SLf\aI.:9�4��aF��\-�R�(�?�#��3����죫��NZ�2��YblVZ:z���j.<�Z�>N�	�g�