XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Ɗ|�݂:�6#�K3�W�&O�]��x�@�2>Ob�,�S�P���	�>M�9���B	I���O����L�(|��w�����FBD��)q@�,�{��U(p6U5M����4�t��ȑ��e�Dq���V��( $�1=��x�O�E��_�ҷq9���2���y[���
���&0�x�K���cMe?�=پS��Q�/�(Ε��%4~�E����t�I�[���?��8�Pm�)<�� �����f�E��,����w<�/���;�⧉�"�U�c�=h��|�e��ﮘ����G^)~��s�d|L�*,�<��r����e`s�އ.�	OZ������m������JQ�ii��m���N�?(�������˩�h�nE�ٚÎ��4��*Ќ�p:�}���-W`�q�7S^̩`�|+/z	�����*���)�|%Hc�#�Y�⫅^}c0:l�[��*�ؽQ]T}�ۈ]�� 6<����W󌙮�	�{��.�}���} ��䊣��Ĝ���! '�3��-	@�/�b�^5?�~sl�E���e��M��؁��}��� ����9nX���qU�D�aҊ���d^��Z�F�/� j6?��Z;���0p{��GMb� |6���Q|���1z?W������w�Q�RU������WN|}4S�#�w2���m=��D$|�`�gp8<�]�1hdo�W�!DgUƁb�b��nĳѤ��I���XlxVHYEB    2327     a90���s7�q �yp���dհ������ށ��jf��*�[����VS���9�H���L����^~�(S���K�yG��wEv0�p������M���xD��|У;��ce�t�Glzj䂘|i��w<���$p/��u�ݢe����)��0�o�8�u���Ź�<|}h����(P�b(M�������v�ɺ. ��R�����IpI�O��!r�P�A��տb�3*:,ձ��Ϋ��2���r;e$��%��È�l!L��W�;JTa��~CĤPk�yO���^X1�
bG��vD�_�4<[}�6�!�����{�7^{�N6���֘kgo�⇍05ƶ��b�RgĚO�'vLyV�K*����dtý�bsU�l��C��6L�"�)�IJ
z��K��������=xf��1�k��B�zp�;��n<D�{q��9pL:���$E���z3��C�� )�b�����#gŁ��"���u%H��A�өG?�H�X��@�su=����
���6O�~|!��`D�9�TPѯ�y+>[�сp����=)�D&��������mAD��y�|n�`��|���� 1RZ�
���zHZ��2@���*?�jO�ͽx_�S��|cC��������:���J�%�/C`1�j�V���[I�_� �aI����xc���"�c:��I��Q����P�=���9.Y��Z� ��iu]2'�_�4Y�[���H�$	��i��;�U,���	Zsc��A%��q�r���'V���o�ԯ���=��_=&�]2	\"�;�}?���%k��.D ���?zF��=v\����b)p��ԍ���?����9��w|�����6]�H����*>�g\���g@x����������)'��1���wl��/;��V�h3Y����A,➁6� �	)Y(����A9��~����&e|� ��Q�N�GcҶ�}��;��k�h�"s�g)L�l��k8�g>����V����t��0iD|���]"i�tw�d��M�NF;x�����3���/\8h0�SS�F&ёU���>�jA��zhM�a��*zL��}��"�O6�@�!�XS�3����A��X��}tĺ�}���}�Ù���_ɖ"����f߅��`�ߺr��9�+���*Y�x��*��yEj��Q��}�]��/$T*��=�K8�i�(}��q.m��p��]�s�L��
\�����)��u/��N��}��[=�_�׬�L5�zOI۬K��6�u�T��irDm�������Ko�H�̈́����t�׳���h({���'��`�R�80%N,�\?*.ˇ��n�&�U��[���Z9�}����az���`�hI=U��`7r�!B�|�#�"M�9YY�W@�hTA�%���?��`��x\����0�}h��1���w��ɓqk��k�y�_6��[��f}�4Ǌ�)�Er�ɀ=���f�nMźyHE�l������(`@|�Ofe:��hG7D�5PP�%���녗1���
��L<~2�����;s7H��\l�?� �Ҍ"g��gN���-E�If�f���E�9��.OR�c��0w���e�l��,{]�P�(��|���ؿ�b��矩	���
�u#u���$�Zcm��,�������~�C^��_ۗ��]>�}���h�ټb���_�`hs��5���.��r��f���s> ��g7�V���"���\q���<�2eukq��:
W�!���tw���OQ�_ԯ9
���gx���1����U��f��E���>A�ݭH���b��x�c���#���/���"���Et�Li�q�H�B�Y���FTt
hL���A"\g�[6����㦵ܙNه3@�C�ߐ��u�?:3���*���b8��e��^�|p�J�L�y�30V������>�c��f���6*�`Zr'�W��B��/ff9�f[��d-�_�e�l��II����>T\xf�K#�J��v�e��.��
jǇ�U�Ao�Jfs��f���8dǇ| r(�!���u�R���h�`4�b���aŔ��fO�,ph_r��M��p�g�� ��Nm��);��y�>����n>,�(	$n'ݲam�O�ԜC���Կ�
�b"����%s�$�	?!����U��6�q\�c.6���G�K�zi#n��O�P�Mm-T��'=ا�]K�M��y��ir����l� �v�H�J�`�wM����z���{w��k�{Y���ՠw(.(�;>1����u�ú��,6bE@�v�L�r�	ϧ��l*M�:�N����u�Ȅ�՜V���χw���bۤtv�F�J��le����K���?4M��d�z̀�5������񟘙��¿�:k���~���@T_y���?���$"j�)����%�D�'$)ڢ���Q�� 9�n�]�]G���i�M?��^(�u�������a
��P;O��=�����W"e�_l��칢�2A`v��!�VK��J ���)��Y��E�j�`��x� �@e䶝�%r@y�����R;U���}�LB����瘎ϯ�(oP���qU�MO�\D���U�MV'���C,F��F��i�$��uu�]1dO�8l��8/r ^yD�����-